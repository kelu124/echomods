// Reading file 'ascii'..

module chip (input io_0_6_1, input io_0_5_1, output io_0_6_0, input io_0_11_1, input io_0_12_0, input io_0_12_1, input io_0_16_0, input io_0_16_1, input io_0_20_0, output io_0_22_0, output io_0_22_1, output io_0_25_1, input io_15_0_1, output io_0_27_1, output io_0_30_0, input io_0_28_1, output io_28_0_0, input io_3_33_1, output io_4_0_1, input io_4_33_0, input io_4_33_1, output io_4_0_0, input io_5_33_0, output io_6_0_1, input io_25_0_0, input io_6_33_0, input io_6_33_1, input io_7_33_0, input io_7_33_1, input io_8_33_0, input io_8_33_1, output io_33_5_0, output io_11_33_1, input io_33_1_1, output io_33_4_1, output io_33_6_0, output io_33_23_1, output io_33_29_1, output io_33_21_1, output io_33_30_0, output io_33_30_1, output io_33_31_0, output io_33_4_0, output io_33_3_1, output io_20_33_1, output io_26_33_0, output io_20_33_0, output io_19_33_1, output io_33_5_1, output io_33_28_0, output io_25_33_0, output io_33_21_0, output io_33_27_1, output io_26_33_1, inout io_27_33_0, inout io_28_33_1, inout io_29_33_0, inout io_29_33_1, output io_30_0_0, inout io_30_33_0, inout io_30_33_1, output io_31_0_0, output io_31_0_1, inout io_31_33_0, inout io_31_33_1, inout io_33_2_1, inout io_33_6_1, inout io_33_10_1, inout io_33_14_1, inout io_33_15_0, inout io_33_15_1, inout io_33_16_0, inout io_33_16_1, output io_33_17_0, output io_33_19_1, output io_33_20_1);

wire n1;
// (0, 0, 'glb_netwk_0')
// (6, 11, 'lutff_global/clk')
// (6, 12, 'lutff_global/clk')
// (7, 8, 'lutff_global/clk')
// (7, 9, 'lutff_global/clk')
// (7, 10, 'lutff_global/clk')
// (7, 11, 'lutff_global/clk')
// (7, 13, 'lutff_global/clk')
// (7, 15, 'lutff_global/clk')
// (9, 12, 'lutff_global/clk')
// (9, 14, 'lutff_global/clk')
// (10, 9, 'lutff_global/clk')
// (10, 10, 'lutff_global/clk')
// (10, 11, 'lutff_global/clk')
// (10, 13, 'lutff_global/clk')
// (10, 14, 'lutff_global/clk')
// (10, 15, 'lutff_global/clk')
// (10, 16, 'lutff_global/clk')
// (10, 17, 'lutff_global/clk')
// (10, 18, 'lutff_global/clk')
// (11, 9, 'lutff_global/clk')
// (11, 10, 'lutff_global/clk')
// (11, 11, 'lutff_global/clk')
// (13, 10, 'lutff_global/clk')
// (14, 10, 'lutff_global/clk')
// (14, 11, 'lutff_global/clk')
// (14, 17, 'lutff_global/clk')
// (15, 10, 'lutff_global/clk')
// (15, 11, 'lutff_global/clk')
// (16, 0, 'span4_horz_r_0')
// (16, 1, 'neigh_op_bnr_0')
// (16, 1, 'neigh_op_bnr_4')
// (16, 8, 'lutff_global/clk')
// (16, 10, 'lutff_global/clk')
// (17, 0, 'fabout')
// (17, 0, 'io_0/D_IN_0')
// (17, 0, 'local_g1_4')
// (17, 0, 'span4_horz_r_4')
// (17, 1, 'neigh_op_bot_0')
// (17, 1, 'neigh_op_bot_4')
// (17, 7, 'lutff_global/clk')
// (17, 9, 'lutff_global/clk')
// (17, 10, 'lutff_global/clk')
// (17, 25, 'lutff_global/clk')
// (18, 0, 'span4_horz_r_8')
// (18, 1, 'neigh_op_bnl_0')
// (18, 1, 'neigh_op_bnl_4')
// (18, 13, 'lutff_global/clk')
// (18, 14, 'lutff_global/clk')
// (18, 16, 'lutff_global/clk')
// (19, 0, 'span4_horz_r_12')
// (19, 8, 'lutff_global/clk')
// (19, 17, 'lutff_global/clk')
// (20, 0, 'span4_horz_l_12')
// (20, 8, 'lutff_global/clk')
// (20, 10, 'lutff_global/clk')
// (20, 14, 'lutff_global/clk')
// (21, 10, 'lutff_global/clk')
// (21, 19, 'lutff_global/clk')
// (22, 10, 'lutff_global/clk')
// (22, 11, 'lutff_global/clk')
// (22, 17, 'lutff_global/clk')
// (22, 18, 'lutff_global/clk')
// (24, 18, 'lutff_global/clk')
// (26, 17, 'lutff_global/clk')

wire n2;
// (0, 0, 'glb_netwk_1')
// (15, 24, 'lutff_global/cen')
// (15, 25, 'lutff_global/cen')
// (15, 26, 'lutff_global/cen')
// (16, 27, 'sp4_r_v_b_46')
// (16, 28, 'sp4_r_v_b_35')
// (16, 29, 'sp4_r_v_b_22')
// (16, 30, 'sp4_r_v_b_11')
// (16, 31, 'sp4_r_v_b_42')
// (16, 32, 'sp4_r_v_b_31')
// (17, 25, 'neigh_op_tnr_0')
// (17, 26, 'neigh_op_rgt_0')
// (17, 26, 'sp4_h_r_5')
// (17, 26, 'sp4_v_t_46')
// (17, 27, 'neigh_op_bnr_0')
// (17, 27, 'sp4_v_b_46')
// (17, 28, 'sp4_v_b_35')
// (17, 29, 'sp4_v_b_22')
// (17, 30, 'sp4_v_b_11')
// (17, 30, 'sp4_v_t_42')
// (17, 31, 'sp4_v_b_42')
// (17, 32, 'sp4_v_b_31')
// (17, 33, 'fabout')
// (17, 33, 'local_g1_2')
// (17, 33, 'span4_vert_18')
// (18, 25, 'neigh_op_top_0')
// (18, 26, 'lutff_0/out')
// (18, 26, 'sp4_h_r_16')
// (18, 27, 'neigh_op_bot_0')
// (19, 25, 'neigh_op_tnl_0')
// (19, 26, 'neigh_op_lft_0')
// (19, 26, 'sp4_h_r_29')
// (19, 27, 'neigh_op_bnl_0')
// (20, 26, 'sp4_h_r_40')
// (21, 26, 'sp4_h_l_40')

wire n3;
// (0, 0, 'glb_netwk_2')
// (5, 17, 'lutff_global/clk')
// (5, 18, 'lutff_global/clk')
// (5, 19, 'lutff_global/clk')
// (7, 16, 'lutff_global/clk')
// (9, 13, 'lutff_global/clk')
// (9, 17, 'lutff_global/clk')
// (9, 18, 'lutff_global/clk')
// (10, 19, 'lutff_global/clk')
// (10, 20, 'lutff_global/clk')
// (10, 23, 'lutff_global/clk')
// (11, 12, 'lutff_global/clk')
// (11, 13, 'lutff_global/clk')
// (11, 16, 'lutff_global/clk')
// (11, 22, 'lutff_global/clk')
// (12, 13, 'lutff_global/clk')
// (12, 17, 'lutff_global/clk')
// (12, 18, 'lutff_global/clk')
// (12, 19, 'lutff_global/clk')
// (12, 20, 'lutff_global/clk')
// (13, 9, 'lutff_global/clk')
// (13, 14, 'lutff_global/clk')
// (13, 15, 'lutff_global/clk')
// (13, 16, 'lutff_global/clk')
// (14, 12, 'lutff_global/clk')
// (14, 13, 'lutff_global/clk')
// (14, 14, 'lutff_global/clk')
// (14, 15, 'lutff_global/clk')
// (14, 16, 'lutff_global/clk')
// (14, 18, 'lutff_global/clk')
// (14, 19, 'lutff_global/clk')
// (14, 20, 'lutff_global/clk')
// (14, 21, 'lutff_global/clk')
// (14, 22, 'lutff_global/clk')
// (14, 23, 'lutff_global/clk')
// (15, 1, 'neigh_op_bnr_2')
// (15, 1, 'neigh_op_bnr_6')
// (15, 9, 'lutff_global/clk')
// (15, 12, 'lutff_global/clk')
// (15, 13, 'lutff_global/clk')
// (15, 14, 'lutff_global/clk')
// (15, 15, 'lutff_global/clk')
// (15, 17, 'lutff_global/clk')
// (15, 18, 'lutff_global/clk')
// (15, 19, 'lutff_global/clk')
// (15, 24, 'lutff_global/clk')
// (15, 25, 'lutff_global/clk')
// (15, 26, 'lutff_global/clk')
// (16, 0, 'io_1/D_IN_0')
// (16, 0, 'span12_vert_12')
// (16, 1, 'neigh_op_bot_2')
// (16, 1, 'neigh_op_bot_6')
// (16, 1, 'sp12_v_b_12')
// (16, 2, 'sp12_v_b_11')
// (16, 3, 'sp12_v_b_8')
// (16, 4, 'sp12_v_b_7')
// (16, 5, 'sp12_v_b_4')
// (16, 6, 'sp12_v_b_3')
// (16, 7, 'sp12_h_r_0')
// (16, 7, 'sp12_v_b_0')
// (16, 9, 'lutff_global/clk')
// (16, 11, 'lutff_global/clk')
// (16, 12, 'lutff_global/clk')
// (16, 13, 'lutff_global/clk')
// (16, 14, 'lutff_global/clk')
// (16, 16, 'lutff_global/clk')
// (16, 17, 'lutff_global/clk')
// (16, 18, 'lutff_global/clk')
// (16, 19, 'lutff_global/clk')
// (16, 20, 'lutff_global/clk')
// (16, 21, 'lutff_global/clk')
// (16, 22, 'lutff_global/clk')
// (16, 23, 'lutff_global/clk')
// (16, 24, 'lutff_global/clk')
// (16, 26, 'lutff_global/clk')
// (17, 1, 'neigh_op_bnl_2')
// (17, 1, 'neigh_op_bnl_6')
// (17, 7, 'sp12_h_r_3')
// (17, 8, 'lutff_global/clk')
// (17, 11, 'lutff_global/clk')
// (17, 12, 'lutff_global/clk')
// (17, 13, 'lutff_global/clk')
// (17, 14, 'lutff_global/clk')
// (17, 15, 'lutff_global/clk')
// (17, 17, 'lutff_global/clk')
// (18, 7, 'lutff_global/clk')
// (18, 7, 'sp12_h_r_4')
// (18, 9, 'lutff_global/clk')
// (18, 11, 'lutff_global/clk')
// (18, 12, 'lutff_global/clk')
// (18, 15, 'lutff_global/clk')
// (18, 17, 'lutff_global/clk')
// (18, 18, 'lutff_global/clk')
// (18, 19, 'lutff_global/clk')
// (18, 20, 'lutff_global/clk')
// (18, 21, 'lutff_global/clk')
// (18, 22, 'lutff_global/clk')
// (18, 23, 'lutff_global/clk')
// (18, 24, 'lutff_global/clk')
// (19, 7, 'sp12_h_r_7')
// (19, 9, 'lutff_global/clk')
// (19, 10, 'lutff_global/clk')
// (19, 11, 'lutff_global/clk')
// (19, 13, 'lutff_global/clk')
// (19, 14, 'lutff_global/clk')
// (19, 15, 'lutff_global/clk')
// (19, 16, 'lutff_global/clk')
// (19, 18, 'lutff_global/clk')
// (19, 19, 'lutff_global/clk')
// (19, 20, 'lutff_global/clk')
// (19, 21, 'lutff_global/clk')
// (19, 22, 'lutff_global/clk')
// (19, 23, 'lutff_global/clk')
// (19, 24, 'lutff_global/clk')
// (19, 25, 'lutff_global/clk')
// (20, 7, 'sp12_h_r_8')
// (20, 11, 'lutff_global/clk')
// (20, 12, 'lutff_global/clk')
// (20, 13, 'lutff_global/clk')
// (20, 16, 'lutff_global/clk')
// (20, 17, 'lutff_global/clk')
// (20, 18, 'lutff_global/clk')
// (20, 19, 'lutff_global/clk')
// (20, 20, 'lutff_global/clk')
// (20, 21, 'lutff_global/clk')
// (20, 22, 'lutff_global/clk')
// (20, 23, 'lutff_global/clk')
// (20, 25, 'lutff_global/clk')
// (20, 26, 'lutff_global/clk')
// (21, 7, 'sp12_h_r_11')
// (21, 11, 'lutff_global/clk')
// (21, 12, 'lutff_global/clk')
// (21, 13, 'lutff_global/clk')
// (21, 14, 'lutff_global/clk')
// (21, 15, 'lutff_global/clk')
// (21, 16, 'lutff_global/clk')
// (21, 17, 'lutff_global/clk')
// (21, 18, 'lutff_global/clk')
// (21, 20, 'lutff_global/clk')
// (21, 21, 'lutff_global/clk')
// (21, 23, 'lutff_global/clk')
// (21, 24, 'lutff_global/clk')
// (22, 7, 'sp12_h_r_12')
// (22, 12, 'lutff_global/clk')
// (22, 13, 'lutff_global/clk')
// (22, 14, 'lutff_global/clk')
// (22, 16, 'lutff_global/clk')
// (22, 19, 'lutff_global/clk')
// (22, 20, 'lutff_global/clk')
// (22, 21, 'lutff_global/clk')
// (22, 22, 'lutff_global/clk')
// (22, 23, 'lutff_global/clk')
// (22, 24, 'lutff_global/clk')
// (23, 7, 'sp12_h_r_15')
// (23, 11, 'lutff_global/clk')
// (23, 12, 'lutff_global/clk')
// (23, 13, 'lutff_global/clk')
// (23, 14, 'lutff_global/clk')
// (23, 15, 'lutff_global/clk')
// (23, 16, 'lutff_global/clk')
// (23, 17, 'lutff_global/clk')
// (23, 18, 'lutff_global/clk')
// (23, 20, 'lutff_global/clk')
// (23, 22, 'lutff_global/clk')
// (24, 7, 'sp12_h_r_16')
// (24, 13, 'lutff_global/clk')
// (24, 14, 'lutff_global/clk')
// (24, 15, 'lutff_global/clk')
// (24, 16, 'lutff_global/clk')
// (24, 17, 'lutff_global/clk')
// (25, 7, 'sp12_h_r_19')
// (26, 7, 'sp12_h_r_20')
// (27, 7, 'sp12_h_r_23')
// (27, 14, 'sp4_r_v_b_39')
// (27, 15, 'sp4_r_v_b_26')
// (27, 16, 'sp4_r_v_b_15')
// (27, 17, 'sp4_r_v_b_2')
// (28, 7, 'sp12_h_l_23')
// (28, 7, 'sp12_v_t_23')
// (28, 8, 'sp12_v_b_23')
// (28, 9, 'sp12_v_b_20')
// (28, 10, 'sp12_v_b_19')
// (28, 11, 'sp12_v_b_16')
// (28, 12, 'sp12_v_b_15')
// (28, 13, 'sp12_v_b_12')
// (28, 13, 'sp4_v_t_39')
// (28, 14, 'sp12_v_b_11')
// (28, 14, 'sp4_v_b_39')
// (28, 15, 'sp12_v_b_8')
// (28, 15, 'sp4_v_b_26')
// (28, 16, 'sp12_v_b_7')
// (28, 16, 'sp4_v_b_15')
// (28, 17, 'sp12_v_b_4')
// (28, 17, 'sp4_h_r_2')
// (28, 17, 'sp4_v_b_2')
// (28, 18, 'sp12_v_b_3')
// (28, 19, 'sp12_v_b_0')
// (29, 17, 'sp4_h_r_15')
// (30, 17, 'sp4_h_r_26')
// (31, 17, 'sp4_h_r_39')
// (32, 17, 'sp4_h_l_39')
// (32, 17, 'sp4_h_r_2')
// (33, 17, 'fabout')
// (33, 17, 'local_g1_2')
// (33, 17, 'span4_horz_2')

wire n4;
// (0, 0, 'glb_netwk_3')
// (0, 17, 'fabout')
// (0, 17, 'local_g1_6')
// (0, 17, 'span4_horz_6')
// (1, 17, 'sp4_h_r_19')
// (2, 17, 'sp4_h_r_30')
// (3, 17, 'sp4_h_r_43')
// (3, 18, 'sp4_r_v_b_37')
// (3, 19, 'sp4_r_v_b_24')
// (3, 20, 'sp4_r_v_b_13')
// (3, 21, 'sp4_r_v_b_0')
// (4, 17, 'sp4_h_l_43')
// (4, 17, 'sp4_v_t_37')
// (4, 18, 'sp4_v_b_37')
// (4, 19, 'sp4_v_b_24')
// (4, 20, 'sp4_v_b_13')
// (4, 21, 'sp12_h_r_1')
// (4, 21, 'sp4_h_r_0')
// (4, 21, 'sp4_v_b_0')
// (5, 17, 'lutff_global/cen')
// (5, 18, 'lutff_global/cen')
// (5, 19, 'lutff_global/cen')
// (5, 21, 'sp12_h_r_2')
// (5, 21, 'sp4_h_r_13')
// (6, 21, 'sp12_h_r_5')
// (6, 21, 'sp4_h_r_24')
// (7, 21, 'sp12_h_r_6')
// (7, 21, 'sp4_h_r_37')
// (8, 21, 'sp12_h_r_9')
// (8, 21, 'sp4_h_l_37')
// (9, 21, 'sp12_h_r_10')
// (10, 21, 'sp12_h_r_13')
// (11, 21, 'sp12_h_r_14')
// (12, 21, 'sp12_h_r_17')
// (13, 21, 'sp12_h_r_18')
// (14, 21, 'sp12_h_r_21')
// (15, 21, 'neigh_op_tnr_3')
// (15, 21, 'sp12_h_r_22')
// (15, 22, 'neigh_op_rgt_3')
// (15, 23, 'neigh_op_bnr_3')
// (16, 21, 'neigh_op_top_3')
// (16, 21, 'sp12_h_l_22')
// (16, 21, 'sp12_v_t_22')
// (16, 22, 'lutff_3/out')
// (16, 22, 'sp12_v_b_22')
// (16, 23, 'neigh_op_bot_3')
// (16, 23, 'sp12_v_b_21')
// (16, 24, 'sp12_v_b_18')
// (16, 25, 'sp12_v_b_17')
// (16, 26, 'sp12_v_b_14')
// (16, 27, 'sp12_v_b_13')
// (16, 28, 'sp12_v_b_10')
// (16, 29, 'sp12_v_b_9')
// (16, 30, 'sp12_v_b_6')
// (16, 31, 'sp12_v_b_5')
// (16, 32, 'sp12_v_b_2')
// (16, 33, 'span12_vert_1')
// (17, 21, 'neigh_op_tnl_3')
// (17, 22, 'neigh_op_lft_3')
// (17, 23, 'neigh_op_bnl_3')

wire n5;
// (0, 0, 'glb_netwk_4')
// (5, 17, 'lutff_global/s_r')
// (5, 18, 'lutff_global/s_r')
// (5, 19, 'lutff_global/s_r')
// (6, 11, 'lutff_global/s_r')
// (6, 12, 'lutff_global/s_r')
// (7, 8, 'lutff_global/s_r')
// (7, 9, 'lutff_global/s_r')
// (7, 10, 'lutff_global/s_r')
// (7, 11, 'lutff_global/s_r')
// (7, 13, 'lutff_global/s_r')
// (7, 15, 'lutff_global/s_r')
// (7, 16, 'lutff_global/s_r')
// (9, 12, 'lutff_global/s_r')
// (9, 13, 'lutff_global/s_r')
// (9, 17, 'lutff_global/s_r')
// (9, 18, 'lutff_global/s_r')
// (10, 9, 'lutff_global/s_r')
// (10, 10, 'lutff_global/s_r')
// (10, 11, 'lutff_global/s_r')
// (10, 13, 'lutff_global/s_r')
// (10, 19, 'lutff_global/s_r')
// (10, 20, 'lutff_global/s_r')
// (10, 23, 'lutff_global/s_r')
// (11, 9, 'lutff_global/s_r')
// (11, 10, 'lutff_global/s_r')
// (11, 11, 'lutff_global/s_r')
// (11, 12, 'lutff_global/s_r')
// (11, 13, 'lutff_global/s_r')
// (11, 16, 'lutff_global/s_r')
// (11, 22, 'lutff_global/s_r')
// (12, 12, 'lutff_global/s_r')
// (12, 13, 'lutff_global/s_r')
// (12, 19, 'lutff_global/s_r')
// (12, 20, 'lutff_global/s_r')
// (13, 9, 'lutff_global/s_r')
// (13, 10, 'lutff_global/s_r')
// (13, 11, 'lutff_global/s_r')
// (13, 12, 'lutff_global/s_r')
// (13, 13, 'lutff_global/s_r')
// (13, 14, 'lutff_global/s_r')
// (13, 16, 'lutff_global/s_r')
// (14, 7, 'lutff_global/s_r')
// (14, 10, 'lutff_global/s_r')
// (14, 11, 'lutff_global/s_r')
// (14, 13, 'lutff_global/s_r')
// (14, 14, 'lutff_global/s_r')
// (14, 16, 'lutff_global/s_r')
// (14, 17, 'lutff_global/s_r')
// (14, 18, 'lutff_global/s_r')
// (14, 19, 'lutff_global/s_r')
// (14, 20, 'lutff_global/s_r')
// (14, 21, 'lutff_global/s_r')
// (14, 22, 'lutff_global/s_r')
// (14, 23, 'lutff_global/s_r')
// (15, 7, 'lutff_global/s_r')
// (15, 9, 'lutff_global/s_r')
// (15, 10, 'lutff_global/s_r')
// (15, 11, 'lutff_global/s_r')
// (15, 12, 'lutff_global/s_r')
// (15, 13, 'lutff_global/s_r')
// (15, 14, 'lutff_global/s_r')
// (15, 15, 'lutff_global/s_r')
// (15, 17, 'lutff_global/s_r')
// (15, 18, 'lutff_global/s_r')
// (15, 19, 'lutff_global/s_r')
// (15, 21, 'neigh_op_tnr_5')
// (15, 22, 'neigh_op_rgt_5')
// (15, 23, 'neigh_op_bnr_5')
// (15, 24, 'lutff_global/s_r')
// (15, 25, 'lutff_global/s_r')
// (15, 26, 'lutff_global/s_r')
// (16, 7, 'lutff_global/s_r')
// (16, 8, 'lutff_global/s_r')
// (16, 9, 'lutff_global/s_r')
// (16, 10, 'lutff_global/s_r')
// (16, 11, 'lutff_global/s_r')
// (16, 12, 'lutff_global/s_r')
// (16, 13, 'lutff_global/s_r')
// (16, 14, 'lutff_global/s_r')
// (16, 15, 'sp12_v_t_22')
// (16, 16, 'lutff_global/s_r')
// (16, 16, 'sp12_v_b_22')
// (16, 17, 'lutff_global/s_r')
// (16, 17, 'sp12_v_b_21')
// (16, 18, 'lutff_global/s_r')
// (16, 18, 'sp12_v_b_18')
// (16, 19, 'lutff_global/s_r')
// (16, 19, 'sp12_v_b_17')
// (16, 20, 'sp12_v_b_14')
// (16, 21, 'lutff_global/s_r')
// (16, 21, 'neigh_op_top_5')
// (16, 21, 'sp12_v_b_13')
// (16, 22, 'lutff_5/out')
// (16, 22, 'sp12_v_b_10')
// (16, 23, 'lutff_global/s_r')
// (16, 23, 'neigh_op_bot_5')
// (16, 23, 'sp12_v_b_9')
// (16, 24, 'lutff_global/s_r')
// (16, 24, 'sp12_v_b_6')
// (16, 25, 'sp12_v_b_5')
// (16, 26, 'lutff_global/s_r')
// (16, 26, 'sp12_v_b_2')
// (16, 27, 'sp12_v_b_1')
// (16, 27, 'sp12_v_t_22')
// (16, 28, 'sp12_v_b_22')
// (16, 29, 'sp12_v_b_21')
// (16, 30, 'sp12_v_b_18')
// (16, 31, 'sp12_v_b_17')
// (16, 32, 'sp12_v_b_14')
// (16, 33, 'fabout')
// (16, 33, 'local_g0_5')
// (16, 33, 'span12_vert_13')
// (17, 7, 'lutff_global/s_r')
// (17, 8, 'lutff_global/s_r')
// (17, 9, 'lutff_global/s_r')
// (17, 10, 'lutff_global/s_r')
// (17, 11, 'lutff_global/s_r')
// (17, 12, 'lutff_global/s_r')
// (17, 13, 'lutff_global/s_r')
// (17, 14, 'lutff_global/s_r')
// (17, 15, 'lutff_global/s_r')
// (17, 17, 'lutff_global/s_r')
// (17, 21, 'neigh_op_tnl_5')
// (17, 22, 'neigh_op_lft_5')
// (17, 23, 'neigh_op_bnl_5')
// (17, 25, 'lutff_global/s_r')
// (18, 7, 'lutff_global/s_r')
// (18, 9, 'lutff_global/s_r')
// (18, 11, 'lutff_global/s_r')
// (18, 12, 'lutff_global/s_r')
// (18, 13, 'lutff_global/s_r')
// (18, 14, 'lutff_global/s_r')
// (18, 15, 'lutff_global/s_r')
// (18, 16, 'lutff_global/s_r')
// (18, 17, 'lutff_global/s_r')
// (18, 18, 'lutff_global/s_r')
// (18, 19, 'lutff_global/s_r')
// (18, 20, 'lutff_global/s_r')
// (18, 22, 'lutff_global/s_r')
// (18, 24, 'lutff_global/s_r')
// (19, 8, 'lutff_global/s_r')
// (19, 9, 'lutff_global/s_r')
// (19, 10, 'lutff_global/s_r')
// (19, 11, 'lutff_global/s_r')
// (19, 13, 'lutff_global/s_r')
// (19, 14, 'lutff_global/s_r')
// (19, 15, 'lutff_global/s_r')
// (19, 16, 'lutff_global/s_r')
// (19, 17, 'lutff_global/s_r')
// (19, 18, 'lutff_global/s_r')
// (19, 19, 'lutff_global/s_r')
// (19, 20, 'lutff_global/s_r')
// (19, 21, 'lutff_global/s_r')
// (19, 22, 'lutff_global/s_r')
// (19, 23, 'lutff_global/s_r')
// (19, 24, 'lutff_global/s_r')
// (19, 25, 'lutff_global/s_r')
// (20, 8, 'lutff_global/s_r')
// (20, 10, 'lutff_global/s_r')
// (20, 11, 'lutff_global/s_r')
// (20, 12, 'lutff_global/s_r')
// (20, 13, 'lutff_global/s_r')
// (20, 14, 'lutff_global/s_r')
// (20, 16, 'lutff_global/s_r')
// (20, 17, 'lutff_global/s_r')
// (20, 18, 'lutff_global/s_r')
// (20, 19, 'lutff_global/s_r')
// (20, 20, 'lutff_global/s_r')
// (20, 21, 'lutff_global/s_r')
// (20, 22, 'lutff_global/s_r')
// (20, 25, 'lutff_global/s_r')
// (20, 26, 'lutff_global/s_r')
// (21, 10, 'lutff_global/s_r')
// (21, 11, 'lutff_global/s_r')
// (21, 12, 'lutff_global/s_r')
// (21, 13, 'lutff_global/s_r')
// (21, 14, 'lutff_global/s_r')
// (21, 15, 'lutff_global/s_r')
// (21, 16, 'lutff_global/s_r')
// (21, 17, 'lutff_global/s_r')
// (21, 18, 'lutff_global/s_r')
// (21, 19, 'lutff_global/s_r')
// (21, 20, 'lutff_global/s_r')
// (21, 21, 'lutff_global/s_r')
// (21, 23, 'lutff_global/s_r')
// (22, 10, 'lutff_global/s_r')
// (22, 11, 'lutff_global/s_r')
// (22, 12, 'lutff_global/s_r')
// (22, 13, 'lutff_global/s_r')
// (22, 14, 'lutff_global/s_r')
// (22, 16, 'lutff_global/s_r')
// (22, 17, 'lutff_global/s_r')
// (22, 18, 'lutff_global/s_r')
// (22, 19, 'lutff_global/s_r')
// (22, 20, 'lutff_global/s_r')
// (22, 21, 'lutff_global/s_r')
// (22, 22, 'lutff_global/s_r')
// (22, 23, 'lutff_global/s_r')
// (22, 24, 'lutff_global/s_r')
// (23, 11, 'lutff_global/s_r')
// (23, 13, 'lutff_global/s_r')
// (23, 14, 'lutff_global/s_r')
// (23, 15, 'lutff_global/s_r')
// (23, 16, 'lutff_global/s_r')
// (23, 17, 'lutff_global/s_r')
// (23, 18, 'lutff_global/s_r')
// (23, 20, 'lutff_global/s_r')
// (23, 22, 'lutff_global/s_r')
// (24, 13, 'lutff_global/s_r')
// (24, 14, 'lutff_global/s_r')
// (24, 15, 'lutff_global/s_r')
// (24, 16, 'lutff_global/s_r')
// (24, 17, 'lutff_global/s_r')
// (24, 18, 'lutff_global/s_r')
// (26, 17, 'lutff_global/s_r')

wire io_0_6_1;
// (0, 0, 'glb_netwk_5')
// (0, 6, 'io_1/D_IN_0')
// (0, 6, 'io_1/PAD')
// (0, 6, 'span12_horz_20')
// (1, 5, 'neigh_op_tnl_2')
// (1, 5, 'neigh_op_tnl_6')
// (1, 6, 'neigh_op_lft_2')
// (1, 6, 'neigh_op_lft_6')
// (1, 6, 'sp12_h_r_23')
// (1, 7, 'neigh_op_bnl_2')
// (1, 7, 'neigh_op_bnl_6')
// (2, 6, 'sp12_h_l_23')
// (2, 6, 'sp12_h_r_0')
// (3, 6, 'sp12_h_r_3')
// (4, 6, 'sp12_h_r_4')
// (5, 6, 'sp12_h_r_7')
// (6, 6, 'sp12_h_r_8')
// (7, 6, 'sp12_h_r_11')
// (8, 6, 'sp12_h_r_12')
// (9, 6, 'sp12_h_r_15')
// (9, 6, 'sp4_h_r_9')
// (10, 6, 'sp12_h_r_16')
// (10, 6, 'sp4_h_r_20')
// (11, 6, 'sp12_h_r_19')
// (11, 6, 'sp4_h_r_33')
// (12, 1, 'sp4_r_v_b_13')
// (12, 2, 'sp4_r_v_b_0')
// (12, 3, 'sp4_r_v_b_44')
// (12, 4, 'sp4_r_v_b_33')
// (12, 5, 'sp4_r_v_b_20')
// (12, 6, 'sp12_h_r_20')
// (12, 6, 'sp4_h_r_44')
// (12, 6, 'sp4_r_v_b_9')
// (12, 12, 'lutff_global/clk')
// (13, 0, 'span4_horz_r_2')
// (13, 0, 'span4_vert_13')
// (13, 1, 'sp4_v_b_13')
// (13, 2, 'sp4_v_b_0')
// (13, 2, 'sp4_v_t_44')
// (13, 3, 'sp4_v_b_44')
// (13, 4, 'sp4_v_b_33')
// (13, 5, 'sp4_v_b_20')
// (13, 6, 'sp12_h_r_23')
// (13, 6, 'sp4_h_l_44')
// (13, 6, 'sp4_v_b_9')
// (13, 11, 'lutff_global/clk')
// (13, 12, 'lutff_global/clk')
// (13, 13, 'lutff_global/clk')
// (14, 0, 'span4_horz_r_6')
// (14, 6, 'sp12_h_l_23')
// (14, 7, 'lutff_global/clk')
// (15, 0, 'span4_horz_r_10')
// (15, 7, 'lutff_global/clk')
// (16, 0, 'fabout')
// (16, 0, 'local_g1_6')
// (16, 0, 'span4_horz_r_14')
// (16, 7, 'lutff_global/clk')
// (17, 0, 'span4_horz_l_14')

wire n7;
// (0, 0, 'glb_netwk_6')
// (0, 16, 'fabout')
// (0, 16, 'local_g0_7')
// (0, 16, 'span4_horz_7')
// (1, 16, 'sp4_h_r_18')
// (2, 16, 'sp4_h_r_31')
// (3, 16, 'sp4_h_r_42')
// (3, 17, 'sp4_r_v_b_42')
// (3, 18, 'sp4_r_v_b_31')
// (3, 19, 'sp4_r_v_b_18')
// (3, 20, 'sp4_r_v_b_7')
// (4, 16, 'sp4_h_l_42')
// (4, 16, 'sp4_v_t_42')
// (4, 17, 'sp4_v_b_42')
// (4, 18, 'sp4_v_b_31')
// (4, 19, 'neigh_op_tnr_1')
// (4, 19, 'sp4_v_b_18')
// (4, 20, 'neigh_op_rgt_1')
// (4, 20, 'sp4_h_r_7')
// (4, 20, 'sp4_v_b_7')
// (4, 21, 'neigh_op_bnr_1')
// (5, 19, 'neigh_op_top_1')
// (5, 20, 'lutff_1/out')
// (5, 20, 'sp4_h_r_18')
// (5, 21, 'neigh_op_bot_1')
// (6, 19, 'neigh_op_tnl_1')
// (6, 20, 'neigh_op_lft_1')
// (6, 20, 'sp4_h_r_31')
// (6, 21, 'neigh_op_bnl_1')
// (7, 20, 'sp4_h_r_42')
// (8, 20, 'sp4_h_l_42')
// (9, 11, 'glb2local_0')
// (9, 11, 'local_g0_4')
// (9, 11, 'lutff_3/in_3')
// (10, 14, 'lutff_global/s_r')
// (10, 15, 'lutff_global/s_r')
// (10, 16, 'lutff_global/s_r')
// (10, 17, 'lutff_global/s_r')
// (10, 18, 'lutff_global/s_r')

wire n8;
// (0, 0, 'glb_netwk_7')
// (14, 17, 'lutff_global/cen')
// (16, 8, 'lutff_global/cen')
// (17, 7, 'lutff_global/cen')
// (17, 10, 'lutff_global/cen')
// (17, 25, 'lutff_global/cen')
// (18, 13, 'lutff_global/cen')
// (18, 14, 'lutff_global/cen')
// (18, 16, 'lutff_global/cen')
// (19, 17, 'lutff_global/cen')
// (20, 8, 'lutff_global/cen')
// (20, 9, 'neigh_op_tnr_1')
// (20, 10, 'neigh_op_rgt_1')
// (20, 11, 'neigh_op_bnr_1')
// (20, 14, 'lutff_global/cen')
// (21, 9, 'neigh_op_top_1')
// (21, 9, 'sp4_r_v_b_46')
// (21, 10, 'lutff_1/out')
// (21, 10, 'sp4_r_v_b_35')
// (21, 11, 'neigh_op_bot_1')
// (21, 11, 'sp4_r_v_b_22')
// (21, 12, 'sp4_r_v_b_11')
// (21, 19, 'lutff_global/cen')
// (22, 8, 'sp4_v_t_46')
// (22, 9, 'neigh_op_tnl_1')
// (22, 9, 'sp4_v_b_46')
// (22, 10, 'neigh_op_lft_1')
// (22, 10, 'sp4_v_b_35')
// (22, 11, 'neigh_op_bnl_1')
// (22, 11, 'sp4_v_b_22')
// (22, 12, 'sp4_h_r_11')
// (22, 12, 'sp4_v_b_11')
// (22, 17, 'lutff_global/cen')
// (22, 18, 'lutff_global/cen')
// (23, 12, 'sp4_h_r_22')
// (24, 12, 'sp4_h_r_35')
// (24, 18, 'lutff_global/cen')
// (25, 12, 'sp4_h_r_46')
// (26, 12, 'sp4_h_l_46')
// (26, 12, 'sp4_h_r_7')
// (26, 17, 'lutff_global/cen')
// (27, 12, 'sp4_h_r_18')
// (28, 12, 'sp4_h_r_31')
// (29, 12, 'sp4_h_r_42')
// (30, 12, 'sp4_h_l_42')
// (30, 12, 'sp4_h_r_7')
// (31, 12, 'sp4_h_r_18')
// (32, 12, 'sp4_h_r_31')
// (33, 12, 'span4_horz_31')
// (33, 12, 'span4_vert_t_13')
// (33, 13, 'span4_vert_b_13')
// (33, 14, 'span4_vert_b_9')
// (33, 15, 'span4_vert_b_5')
// (33, 16, 'fabout')
// (33, 16, 'local_g0_1')
// (33, 16, 'span4_vert_b_1')

wire io_0_5_1;
// (0, 5, 'io_1/D_IN_0')
// (0, 5, 'io_1/PAD')
// (0, 5, 'span12_horz_20')
// (1, 4, 'neigh_op_tnl_2')
// (1, 4, 'neigh_op_tnl_6')
// (1, 5, 'neigh_op_lft_2')
// (1, 5, 'neigh_op_lft_6')
// (1, 5, 'sp12_h_r_23')
// (1, 6, 'neigh_op_bnl_2')
// (1, 6, 'neigh_op_bnl_6')
// (2, 5, 'sp12_h_l_23')
// (2, 5, 'sp12_h_r_0')
// (3, 5, 'sp12_h_r_3')
// (4, 5, 'sp12_h_r_4')
// (5, 5, 'sp12_h_r_7')
// (6, 5, 'sp12_h_r_8')
// (7, 5, 'sp12_h_r_11')
// (8, 5, 'sp12_h_r_12')
// (9, 5, 'sp12_h_r_15')
// (9, 5, 'sp4_h_r_9')
// (10, 5, 'sp12_h_r_16')
// (10, 5, 'sp4_h_r_20')
// (11, 5, 'sp12_h_r_19')
// (11, 5, 'sp4_h_r_33')
// (12, 5, 'sp12_h_r_20')
// (12, 5, 'sp4_h_r_44')
// (12, 6, 'sp4_r_v_b_39')
// (12, 7, 'sp4_r_v_b_26')
// (12, 8, 'sp4_r_v_b_15')
// (12, 9, 'sp4_r_v_b_2')
// (12, 10, 'sp4_r_v_b_47')
// (12, 11, 'sp4_r_v_b_34')
// (12, 12, 'local_g3_7')
// (12, 12, 'lutff_3/in_3')
// (12, 12, 'sp4_r_v_b_23')
// (12, 13, 'sp4_r_v_b_10')
// (13, 5, 'sp12_h_r_23')
// (13, 5, 'sp4_h_l_44')
// (13, 5, 'sp4_v_t_39')
// (13, 6, 'sp4_v_b_39')
// (13, 7, 'sp4_v_b_26')
// (13, 8, 'sp4_v_b_15')
// (13, 9, 'sp4_v_b_2')
// (13, 9, 'sp4_v_t_47')
// (13, 10, 'sp4_v_b_47')
// (13, 11, 'sp4_v_b_34')
// (13, 12, 'sp4_v_b_23')
// (13, 13, 'sp4_v_b_10')
// (14, 5, 'sp12_h_l_23')

wire io_0_6_0;
// (0, 6, 'io_0/D_OUT_0')
// (0, 6, 'io_0/PAD')
// (0, 6, 'local_g0_6')
// (0, 6, 'span12_horz_22')
// (1, 6, 'sp12_h_l_22')
// (1, 6, 'sp12_h_r_1')
// (2, 6, 'sp12_h_r_2')
// (3, 6, 'sp12_h_r_5')
// (4, 6, 'sp12_h_r_6')
// (5, 6, 'sp12_h_r_9')
// (6, 6, 'sp12_h_r_10')
// (6, 7, 'sp12_h_r_1')
// (6, 7, 'sp12_v_t_22')
// (6, 8, 'local_g2_6')
// (6, 8, 'lutff_1/in_3')
// (6, 8, 'sp12_v_b_22')
// (6, 9, 'sp12_v_b_21')
// (6, 10, 'sp12_v_b_18')
// (6, 11, 'sp12_v_b_17')
// (6, 12, 'sp12_v_b_14')
// (6, 13, 'sp12_v_b_13')
// (6, 14, 'sp12_v_b_10')
// (6, 15, 'sp12_v_b_9')
// (6, 16, 'sp12_v_b_6')
// (6, 17, 'sp12_v_b_5')
// (6, 18, 'sp12_v_b_2')
// (6, 19, 'sp12_v_b_1')
// (7, 6, 'sp12_h_r_13')
// (7, 7, 'sp12_h_r_2')
// (8, 6, 'sp12_h_r_14')
// (8, 7, 'sp12_h_r_5')
// (9, 6, 'sp12_h_r_17')
// (9, 7, 'sp12_h_r_6')
// (10, 6, 'sp12_h_r_18')
// (10, 7, 'sp12_h_r_9')
// (11, 6, 'sp12_h_r_21')
// (11, 7, 'sp12_h_r_10')
// (12, 6, 'neigh_op_tnr_3')
// (12, 6, 'sp12_h_r_22')
// (12, 7, 'neigh_op_rgt_3')
// (12, 7, 'sp12_h_r_13')
// (12, 8, 'neigh_op_bnr_3')
// (13, 6, 'neigh_op_top_3')
// (13, 6, 'sp12_h_l_22')
// (13, 6, 'sp12_v_t_22')
// (13, 7, 'lutff_3/out')
// (13, 7, 'sp12_h_r_14')
// (13, 7, 'sp12_v_b_22')
// (13, 8, 'neigh_op_bot_3')
// (13, 8, 'sp12_v_b_21')
// (13, 9, 'sp12_v_b_18')
// (13, 10, 'sp12_v_b_17')
// (13, 11, 'sp12_v_b_14')
// (13, 12, 'sp12_v_b_13')
// (13, 13, 'sp12_v_b_10')
// (13, 14, 'sp12_v_b_9')
// (13, 15, 'sp12_v_b_6')
// (13, 16, 'sp12_v_b_5')
// (13, 17, 'sp12_v_b_2')
// (13, 18, 'sp12_v_b_1')
// (14, 6, 'neigh_op_tnl_3')
// (14, 7, 'neigh_op_lft_3')
// (14, 7, 'sp12_h_r_17')
// (14, 8, 'neigh_op_bnl_3')
// (15, 7, 'sp12_h_r_18')
// (16, 7, 'sp12_h_r_21')
// (17, 7, 'sp12_h_r_22')
// (18, 7, 'sp12_h_l_22')

wire io_0_11_1;
// (0, 11, 'io_1/D_IN_0')
// (0, 11, 'io_1/PAD')
// (0, 11, 'span12_horz_12')
// (1, 10, 'neigh_op_tnl_2')
// (1, 10, 'neigh_op_tnl_6')
// (1, 11, 'neigh_op_lft_2')
// (1, 11, 'neigh_op_lft_6')
// (1, 11, 'sp12_h_r_15')
// (1, 12, 'neigh_op_bnl_2')
// (1, 12, 'neigh_op_bnl_6')
// (2, 11, 'sp12_h_r_16')
// (3, 11, 'sp12_h_r_19')
// (4, 11, 'sp12_h_r_20')
// (5, 11, 'sp12_h_r_23')
// (6, 11, 'sp12_h_l_23')
// (6, 11, 'sp12_v_t_23')
// (6, 12, 'sp12_v_b_23')
// (6, 13, 'sp12_v_b_20')
// (6, 14, 'sp12_v_b_19')
// (6, 15, 'sp12_v_b_16')
// (6, 16, 'sp12_v_b_15')
// (6, 17, 'sp12_v_b_12')
// (6, 18, 'sp12_v_b_11')
// (6, 19, 'sp12_v_b_8')
// (6, 20, 'sp12_v_b_7')
// (6, 21, 'sp12_v_b_4')
// (6, 22, 'sp12_v_b_3')
// (6, 23, 'sp12_h_r_0')
// (6, 23, 'sp12_v_b_0')
// (7, 23, 'sp12_h_r_3')
// (8, 23, 'sp12_h_r_4')
// (9, 23, 'sp12_h_r_7')
// (10, 23, 'sp12_h_r_8')
// (11, 23, 'sp12_h_r_11')
// (12, 23, 'sp12_h_r_12')
// (13, 23, 'sp12_h_r_15')
// (14, 23, 'sp12_h_r_16')
// (15, 23, 'sp12_h_r_19')
// (16, 23, 'local_g1_4')
// (16, 23, 'lutff_4/in_3')
// (16, 23, 'sp12_h_r_20')
// (17, 23, 'sp12_h_r_23')
// (18, 23, 'sp12_h_l_23')

wire io_0_12_0;
// (0, 12, 'io_0/D_IN_0')
// (0, 12, 'io_0/PAD')
// (0, 12, 'span12_horz_16')
// (1, 11, 'neigh_op_tnl_0')
// (1, 11, 'neigh_op_tnl_4')
// (1, 12, 'neigh_op_lft_0')
// (1, 12, 'neigh_op_lft_4')
// (1, 12, 'sp12_h_r_19')
// (1, 13, 'neigh_op_bnl_0')
// (1, 13, 'neigh_op_bnl_4')
// (2, 12, 'sp12_h_r_20')
// (3, 12, 'sp12_h_r_23')
// (4, 12, 'sp12_h_l_23')
// (4, 12, 'sp12_v_t_23')
// (4, 13, 'sp12_v_b_23')
// (4, 14, 'sp12_v_b_20')
// (4, 15, 'sp12_v_b_19')
// (4, 16, 'sp12_v_b_16')
// (4, 17, 'sp12_v_b_15')
// (4, 18, 'sp12_v_b_12')
// (4, 19, 'sp12_v_b_11')
// (4, 20, 'sp12_v_b_8')
// (4, 21, 'sp12_v_b_7')
// (4, 22, 'sp12_v_b_4')
// (4, 23, 'sp12_v_b_3')
// (4, 24, 'sp12_h_r_0')
// (4, 24, 'sp12_v_b_0')
// (5, 24, 'sp12_h_r_3')
// (6, 24, 'sp12_h_r_4')
// (7, 24, 'sp12_h_r_7')
// (8, 24, 'sp12_h_r_8')
// (9, 24, 'sp12_h_r_11')
// (10, 24, 'sp12_h_r_12')
// (11, 24, 'sp12_h_r_15')
// (12, 24, 'sp12_h_r_16')
// (13, 24, 'sp12_h_r_19')
// (13, 24, 'sp4_h_r_11')
// (14, 24, 'sp12_h_r_20')
// (14, 24, 'sp4_h_r_22')
// (15, 24, 'sp12_h_r_23')
// (15, 24, 'sp4_h_r_35')
// (16, 21, 'sp4_r_v_b_46')
// (16, 22, 'sp4_r_v_b_35')
// (16, 23, 'local_g3_6')
// (16, 23, 'lutff_3/in_0')
// (16, 23, 'sp4_r_v_b_22')
// (16, 24, 'sp12_h_l_23')
// (16, 24, 'sp4_h_r_46')
// (16, 24, 'sp4_r_v_b_11')
// (17, 20, 'sp4_v_t_46')
// (17, 21, 'sp4_v_b_46')
// (17, 22, 'sp4_v_b_35')
// (17, 23, 'sp4_v_b_22')
// (17, 24, 'sp4_h_l_46')
// (17, 24, 'sp4_v_b_11')

wire io_0_12_1;
// (0, 12, 'io_1/D_IN_0')
// (0, 12, 'io_1/PAD')
// (0, 12, 'span12_horz_12')
// (1, 11, 'neigh_op_tnl_2')
// (1, 11, 'neigh_op_tnl_6')
// (1, 12, 'neigh_op_lft_2')
// (1, 12, 'neigh_op_lft_6')
// (1, 12, 'sp12_h_r_15')
// (1, 13, 'neigh_op_bnl_2')
// (1, 13, 'neigh_op_bnl_6')
// (2, 12, 'sp12_h_r_16')
// (3, 12, 'sp12_h_r_19')
// (4, 12, 'sp12_h_r_20')
// (5, 12, 'sp12_h_r_23')
// (6, 0, 'span12_vert_23')
// (6, 1, 'sp12_v_b_23')
// (6, 2, 'sp12_v_b_20')
// (6, 3, 'sp12_v_b_19')
// (6, 4, 'sp12_v_b_16')
// (6, 5, 'sp12_v_b_15')
// (6, 6, 'sp12_v_b_12')
// (6, 7, 'sp12_v_b_11')
// (6, 8, 'local_g3_0')
// (6, 8, 'lutff_1/in_0')
// (6, 8, 'sp12_v_b_8')
// (6, 9, 'sp12_v_b_7')
// (6, 10, 'sp12_v_b_4')
// (6, 11, 'sp12_v_b_3')
// (6, 12, 'sp12_h_l_23')
// (6, 12, 'sp12_v_b_0')

reg n14 = 0;
// (0, 12, 'span12_horz_1')
// (1, 12, 'sp12_h_r_2')
// (2, 12, 'sp12_h_r_5')
// (3, 12, 'sp12_h_r_6')
// (4, 12, 'sp12_h_r_9')
// (5, 12, 'sp12_h_r_10')
// (6, 12, 'sp12_h_r_13')
// (7, 12, 'local_g0_6')
// (7, 12, 'lutff_1/in_3')
// (7, 12, 'sp12_h_r_14')
// (8, 12, 'sp12_h_r_17')
// (9, 12, 'sp12_h_r_18')
// (10, 12, 'sp12_h_r_21')
// (11, 9, 'sp4_h_r_9')
// (11, 12, 'sp12_h_r_22')
// (11, 13, 'sp4_h_r_8')
// (12, 9, 'sp4_h_r_20')
// (12, 12, 'sp12_h_l_22')
// (12, 12, 'sp12_h_r_1')
// (12, 13, 'sp4_h_r_21')
// (13, 9, 'local_g2_1')
// (13, 9, 'lutff_0/in_3')
// (13, 9, 'sp4_h_r_33')
// (13, 12, 'sp12_h_r_2')
// (13, 13, 'local_g3_0')
// (13, 13, 'lutff_2/in_3')
// (13, 13, 'sp4_h_r_32')
// (14, 9, 'sp4_h_r_44')
// (14, 10, 'sp4_r_v_b_38')
// (14, 11, 'neigh_op_tnr_7')
// (14, 11, 'sp4_r_v_b_27')
// (14, 12, 'neigh_op_rgt_7')
// (14, 12, 'sp12_h_r_5')
// (14, 12, 'sp4_r_v_b_14')
// (14, 13, 'neigh_op_bnr_7')
// (14, 13, 'sp4_h_r_45')
// (14, 13, 'sp4_r_v_b_3')
// (15, 9, 'sp4_h_l_44')
// (15, 9, 'sp4_v_t_38')
// (15, 10, 'sp4_v_b_38')
// (15, 11, 'neigh_op_top_7')
// (15, 11, 'sp4_v_b_27')
// (15, 12, 'lutff_7/out')
// (15, 12, 'sp12_h_r_6')
// (15, 12, 'sp4_v_b_14')
// (15, 13, 'neigh_op_bot_7')
// (15, 13, 'sp4_h_l_45')
// (15, 13, 'sp4_v_b_3')
// (16, 11, 'neigh_op_tnl_7')
// (16, 12, 'neigh_op_lft_7')
// (16, 12, 'sp12_h_r_9')
// (16, 13, 'neigh_op_bnl_7')
// (17, 12, 'sp12_h_r_10')
// (18, 12, 'sp12_h_r_13')
// (19, 12, 'sp12_h_r_14')
// (20, 12, 'sp12_h_r_17')
// (21, 12, 'sp12_h_r_18')
// (22, 12, 'sp12_h_r_21')
// (23, 12, 'sp12_h_r_22')
// (24, 12, 'sp12_h_l_22')

wire io_0_16_0;
// (0, 16, 'io_0/D_IN_0')
// (0, 16, 'io_0/PAD')
// (0, 16, 'span12_horz_0')
// (1, 15, 'neigh_op_tnl_0')
// (1, 15, 'neigh_op_tnl_4')
// (1, 16, 'neigh_op_lft_0')
// (1, 16, 'neigh_op_lft_4')
// (1, 16, 'sp12_h_r_3')
// (1, 17, 'neigh_op_bnl_0')
// (1, 17, 'neigh_op_bnl_4')
// (2, 16, 'sp12_h_r_4')
// (3, 16, 'sp12_h_r_7')
// (4, 16, 'sp12_h_r_8')
// (5, 16, 'sp12_h_r_11')
// (6, 16, 'local_g1_4')
// (6, 16, 'lutff_0/in_1')
// (6, 16, 'sp12_h_r_12')
// (7, 16, 'local_g0_7')
// (7, 16, 'lutff_7/in_0')
// (7, 16, 'sp12_h_r_15')
// (8, 16, 'sp12_h_r_16')
// (9, 16, 'local_g0_3')
// (9, 16, 'local_g1_3')
// (9, 16, 'lutff_3/in_1')
// (9, 16, 'lutff_4/in_1')
// (9, 16, 'sp12_h_r_19')
// (10, 16, 'sp12_h_r_20')
// (11, 16, 'sp12_h_r_23')
// (12, 16, 'sp12_h_l_23')

wire io_0_16_1;
// (0, 16, 'io_1/D_IN_0')
// (0, 16, 'io_1/PAD')
// (0, 16, 'span12_horz_20')
// (1, 15, 'neigh_op_tnl_2')
// (1, 15, 'neigh_op_tnl_6')
// (1, 16, 'neigh_op_lft_2')
// (1, 16, 'neigh_op_lft_6')
// (1, 16, 'sp12_h_r_23')
// (1, 17, 'neigh_op_bnl_2')
// (1, 17, 'neigh_op_bnl_6')
// (2, 4, 'sp12_h_r_0')
// (2, 4, 'sp12_v_t_23')
// (2, 5, 'sp12_v_b_23')
// (2, 6, 'sp12_v_b_20')
// (2, 7, 'sp12_v_b_19')
// (2, 8, 'sp12_v_b_16')
// (2, 9, 'sp12_v_b_15')
// (2, 10, 'sp12_v_b_12')
// (2, 11, 'sp12_v_b_11')
// (2, 12, 'sp12_v_b_8')
// (2, 13, 'sp12_v_b_7')
// (2, 14, 'sp12_v_b_4')
// (2, 15, 'sp12_v_b_3')
// (2, 16, 'sp12_h_l_23')
// (2, 16, 'sp12_v_b_0')
// (3, 4, 'sp12_h_r_3')
// (4, 4, 'sp12_h_r_4')
// (5, 4, 'sp12_h_r_7')
// (6, 4, 'sp12_h_r_8')
// (7, 4, 'sp12_h_r_11')
// (8, 4, 'sp12_h_r_12')
// (9, 4, 'sp12_h_r_15')
// (9, 4, 'sp4_h_r_9')
// (10, 4, 'sp12_h_r_16')
// (10, 4, 'sp4_h_r_20')
// (11, 4, 'sp12_h_r_19')
// (11, 4, 'sp4_h_r_33')
// (12, 1, 'sp4_r_v_b_38')
// (12, 2, 'sp4_r_v_b_27')
// (12, 3, 'sp4_r_v_b_14')
// (12, 4, 'sp12_h_r_20')
// (12, 4, 'sp4_h_r_44')
// (12, 4, 'sp4_r_v_b_3')
// (13, 0, 'fabout')
// (13, 0, 'local_g1_6')
// (13, 0, 'span4_vert_38')
// (13, 1, 'sp4_v_b_38')
// (13, 2, 'sp4_v_b_27')
// (13, 3, 'sp4_v_b_14')
// (13, 4, 'sp12_h_r_23')
// (13, 4, 'sp4_h_l_44')
// (13, 4, 'sp4_v_b_3')
// (14, 4, 'sp12_h_l_23')

reg n17 = 0;
// (0, 17, 'span12_horz_3')
// (1, 17, 'sp12_h_r_4')
// (2, 17, 'sp12_h_r_7')
// (3, 17, 'sp12_h_r_8')
// (4, 16, 'neigh_op_tnr_2')
// (4, 17, 'neigh_op_rgt_2')
// (4, 17, 'sp12_h_r_11')
// (4, 18, 'neigh_op_bnr_2')
// (5, 16, 'neigh_op_top_2')
// (5, 17, 'local_g1_2')
// (5, 17, 'lutff_2/in_1')
// (5, 17, 'lutff_2/out')
// (5, 17, 'sp12_h_r_12')
// (5, 18, 'neigh_op_bot_2')
// (6, 16, 'neigh_op_tnl_2')
// (6, 17, 'neigh_op_lft_2')
// (6, 17, 'sp12_h_r_15')
// (6, 18, 'neigh_op_bnl_2')
// (7, 17, 'sp12_h_r_16')
// (8, 17, 'sp12_h_r_19')
// (9, 17, 'sp12_h_r_20')
// (10, 17, 'sp12_h_r_23')
// (11, 17, 'sp12_h_l_23')
// (11, 17, 'sp12_h_r_0')
// (12, 17, 'sp12_h_r_3')
// (13, 17, 'sp12_h_r_4')
// (14, 17, 'sp12_h_r_7')
// (14, 17, 'sp4_h_r_5')
// (15, 17, 'sp12_h_r_8')
// (15, 17, 'sp4_h_r_16')
// (16, 17, 'sp12_h_r_11')
// (16, 17, 'sp4_h_r_29')
// (17, 17, 'sp12_h_r_12')
// (17, 17, 'sp4_h_r_40')
// (17, 18, 'sp4_r_v_b_40')
// (17, 19, 'sp4_r_v_b_29')
// (17, 20, 'sp4_r_v_b_16')
// (17, 21, 'sp4_r_v_b_5')
// (18, 17, 'sp12_h_r_15')
// (18, 17, 'sp4_h_l_40')
// (18, 17, 'sp4_v_t_40')
// (18, 18, 'sp4_v_b_40')
// (18, 19, 'sp4_v_b_29')
// (18, 20, 'sp4_v_b_16')
// (18, 21, 'local_g1_5')
// (18, 21, 'lutff_3/in_3')
// (18, 21, 'sp4_v_b_5')
// (19, 17, 'sp12_h_r_16')
// (20, 17, 'sp12_h_r_19')
// (21, 17, 'sp12_h_r_20')
// (22, 17, 'sp12_h_r_23')
// (23, 17, 'sp12_h_l_23')

wire io_0_20_0;
// (0, 20, 'io_0/D_IN_0')
// (0, 20, 'io_0/PAD')
// (0, 20, 'span4_horz_16')
// (1, 19, 'neigh_op_tnl_0')
// (1, 19, 'neigh_op_tnl_4')
// (1, 20, 'neigh_op_lft_0')
// (1, 20, 'neigh_op_lft_4')
// (1, 20, 'sp4_h_r_29')
// (1, 21, 'neigh_op_bnl_0')
// (1, 21, 'neigh_op_bnl_4')
// (2, 17, 'sp4_r_v_b_46')
// (2, 18, 'sp4_r_v_b_35')
// (2, 19, 'sp4_r_v_b_22')
// (2, 20, 'sp4_h_r_40')
// (2, 20, 'sp4_r_v_b_11')
// (3, 16, 'sp4_h_r_11')
// (3, 16, 'sp4_v_t_46')
// (3, 17, 'sp4_v_b_46')
// (3, 18, 'sp4_v_b_35')
// (3, 19, 'sp4_v_b_22')
// (3, 20, 'sp4_h_l_40')
// (3, 20, 'sp4_v_b_11')
// (4, 16, 'sp4_h_r_22')
// (5, 16, 'sp4_h_r_35')
// (6, 16, 'local_g3_6')
// (6, 16, 'lutff_0/in_3')
// (6, 16, 'sp4_h_r_46')
// (7, 16, 'local_g1_7')
// (7, 16, 'lutff_7/in_3')
// (7, 16, 'sp4_h_l_46')
// (7, 16, 'sp4_h_r_7')
// (8, 16, 'sp4_h_r_18')
// (9, 16, 'local_g2_7')
// (9, 16, 'lutff_3/in_0')
// (9, 16, 'lutff_4/in_3')
// (9, 16, 'sp4_h_r_31')
// (10, 16, 'sp4_h_r_42')
// (11, 16, 'sp4_h_l_42')

wire io_0_22_0;
// (0, 21, 'span4_horz_1')
// (0, 21, 'span4_vert_t_12')
// (0, 22, 'io_0/D_OUT_0')
// (0, 22, 'io_0/PAD')
// (0, 22, 'local_g0_4')
// (0, 22, 'span4_vert_b_12')
// (0, 23, 'span4_vert_b_8')
// (0, 24, 'span4_vert_b_4')
// (0, 25, 'span4_vert_b_0')
// (1, 21, 'sp12_h_r_0')
// (1, 21, 'sp4_h_r_12')
// (2, 21, 'sp12_h_r_3')
// (2, 21, 'sp4_h_r_25')
// (3, 21, 'sp12_h_r_4')
// (3, 21, 'sp4_h_r_36')
// (4, 21, 'sp12_h_r_7')
// (4, 21, 'sp4_h_l_36')
// (5, 21, 'sp12_h_r_8')
// (6, 21, 'sp12_h_r_11')
// (7, 21, 'sp12_h_r_12')
// (8, 21, 'sp12_h_r_15')
// (9, 21, 'sp12_h_r_16')
// (10, 21, 'sp12_h_r_19')
// (11, 21, 'sp12_h_r_20')
// (12, 20, 'neigh_op_tnr_0')
// (12, 21, 'neigh_op_rgt_0')
// (12, 21, 'sp12_h_r_23')
// (12, 22, 'neigh_op_bnr_0')
// (13, 9, 'sp12_v_t_23')
// (13, 10, 'sp12_v_b_23')
// (13, 11, 'sp12_v_b_20')
// (13, 12, 'sp12_v_b_19')
// (13, 13, 'sp12_v_b_16')
// (13, 14, 'sp12_v_b_15')
// (13, 15, 'sp12_v_b_12')
// (13, 16, 'sp12_v_b_11')
// (13, 17, 'sp12_v_b_8')
// (13, 18, 'sp12_v_b_7')
// (13, 19, 'sp12_v_b_4')
// (13, 20, 'neigh_op_top_0')
// (13, 20, 'sp12_v_b_3')
// (13, 21, 'lutff_0/out')
// (13, 21, 'sp12_h_l_23')
// (13, 21, 'sp12_v_b_0')
// (13, 22, 'neigh_op_bot_0')
// (14, 20, 'neigh_op_tnl_0')
// (14, 21, 'neigh_op_lft_0')
// (14, 22, 'neigh_op_bnl_0')

wire io_0_22_1;
// (0, 21, 'span4_vert_t_13')
// (0, 22, 'io_1/D_OUT_0')
// (0, 22, 'io_1/PAD')
// (0, 22, 'local_g0_5')
// (0, 22, 'span4_vert_b_13')
// (0, 23, 'span4_vert_b_9')
// (0, 24, 'span4_vert_b_5')
// (0, 25, 'span4_horz_7')
// (0, 25, 'span4_vert_b_1')
// (1, 25, 'sp4_h_r_18')
// (2, 25, 'sp4_h_r_31')
// (3, 25, 'sp4_h_r_42')
// (4, 25, 'sp4_h_l_42')
// (4, 25, 'sp4_h_r_11')
// (5, 25, 'sp4_h_r_22')
// (6, 25, 'sp4_h_r_35')
// (7, 25, 'sp4_h_r_46')
// (8, 25, 'sp4_h_l_46')
// (8, 25, 'sp4_h_r_8')
// (9, 25, 'sp4_h_r_21')
// (10, 25, 'sp4_h_r_32')
// (11, 25, 'sp4_h_r_45')
// (12, 24, 'neigh_op_tnr_0')
// (12, 25, 'neigh_op_rgt_0')
// (12, 25, 'sp4_h_l_45')
// (12, 25, 'sp4_h_r_5')
// (12, 26, 'neigh_op_bnr_0')
// (13, 24, 'neigh_op_top_0')
// (13, 25, 'lutff_0/out')
// (13, 25, 'sp4_h_r_16')
// (13, 26, 'neigh_op_bot_0')
// (14, 24, 'neigh_op_tnl_0')
// (14, 25, 'neigh_op_lft_0')
// (14, 25, 'sp4_h_r_29')
// (14, 26, 'neigh_op_bnl_0')
// (15, 25, 'sp4_h_r_40')
// (16, 25, 'sp4_h_l_40')

wire io_0_25_1;
assign io_0_25_1 = io_15_0_1;
// (0, 23, 'span4_horz_25')
// (0, 23, 'span4_vert_t_12')
// (0, 24, 'span4_vert_b_12')
// (0, 25, 'io_1/D_OUT_0')
// (0, 25, 'io_1/PAD')
// (0, 25, 'local_g1_0')
// (0, 25, 'span4_vert_b_8')
// (0, 26, 'span4_vert_b_4')
// (0, 27, 'span4_vert_b_0')
// (1, 23, 'sp4_h_r_36')
// (2, 23, 'sp4_h_l_36')
// (2, 23, 'sp4_h_r_5')
// (3, 11, 'sp12_h_r_0')
// (3, 23, 'sp4_h_r_16')
// (4, 11, 'sp12_h_r_3')
// (4, 23, 'sp4_h_r_29')
// (5, 11, 'sp12_h_r_4')
// (5, 20, 'local_g3_0')
// (5, 20, 'lutff_1/in_0')
// (5, 20, 'sp4_r_v_b_40')
// (5, 21, 'sp4_r_v_b_29')
// (5, 22, 'sp4_r_v_b_16')
// (5, 23, 'sp4_h_r_40')
// (5, 23, 'sp4_r_v_b_5')
// (6, 11, 'sp12_h_r_7')
// (6, 19, 'sp4_h_r_5')
// (6, 19, 'sp4_v_t_40')
// (6, 20, 'sp4_v_b_40')
// (6, 21, 'sp4_v_b_29')
// (6, 22, 'sp4_v_b_16')
// (6, 23, 'sp4_h_l_40')
// (6, 23, 'sp4_v_b_5')
// (7, 11, 'sp12_h_r_8')
// (7, 19, 'sp4_h_r_11')
// (7, 19, 'sp4_h_r_16')
// (8, 11, 'sp12_h_r_11')
// (8, 19, 'sp4_h_r_22')
// (8, 19, 'sp4_h_r_29')
// (9, 11, 'local_g1_4')
// (9, 11, 'lutff_3/in_0')
// (9, 11, 'sp12_h_r_12')
// (9, 19, 'local_g2_3')
// (9, 19, 'lutff_2/in_1')
// (9, 19, 'sp4_h_r_35')
// (9, 19, 'sp4_h_r_40')
// (10, 11, 'sp12_h_r_15')
// (10, 12, 'sp4_r_v_b_37')
// (10, 12, 'sp4_r_v_b_43')
// (10, 13, 'sp4_r_v_b_24')
// (10, 13, 'sp4_r_v_b_30')
// (10, 14, 'local_g3_3')
// (10, 14, 'lutff_1/in_1')
// (10, 14, 'lutff_2/in_2')
// (10, 14, 'lutff_3/in_3')
// (10, 14, 'sp4_r_v_b_13')
// (10, 14, 'sp4_r_v_b_19')
// (10, 15, 'local_g0_6')
// (10, 15, 'local_g1_0')
// (10, 15, 'lutff_0/in_3')
// (10, 15, 'lutff_1/in_0')
// (10, 15, 'lutff_2/in_0')
// (10, 15, 'lutff_3/in_0')
// (10, 15, 'lutff_4/in_0')
// (10, 15, 'lutff_5/in_0')
// (10, 15, 'lutff_6/in_0')
// (10, 15, 'lutff_7/in_0')
// (10, 15, 'sp4_h_r_6')
// (10, 15, 'sp4_r_v_b_0')
// (10, 15, 'sp4_r_v_b_6')
// (10, 16, 'local_g2_7')
// (10, 16, 'local_g3_3')
// (10, 16, 'lutff_0/in_0')
// (10, 16, 'lutff_1/in_0')
// (10, 16, 'lutff_2/in_0')
// (10, 16, 'lutff_3/in_0')
// (10, 16, 'lutff_4/in_0')
// (10, 16, 'lutff_5/in_0')
// (10, 16, 'lutff_6/in_0')
// (10, 16, 'lutff_7/in_0')
// (10, 16, 'sp4_r_v_b_39')
// (10, 16, 'sp4_r_v_b_43')
// (10, 17, 'local_g0_2')
// (10, 17, 'local_g1_6')
// (10, 17, 'lutff_0/in_0')
// (10, 17, 'lutff_1/in_0')
// (10, 17, 'lutff_2/in_0')
// (10, 17, 'lutff_3/in_0')
// (10, 17, 'lutff_4/in_0')
// (10, 17, 'lutff_5/in_0')
// (10, 17, 'sp4_r_v_b_26')
// (10, 17, 'sp4_r_v_b_30')
// (10, 18, 'sp4_r_v_b_15')
// (10, 18, 'sp4_r_v_b_19')
// (10, 19, 'sp4_h_l_40')
// (10, 19, 'sp4_h_r_2')
// (10, 19, 'sp4_h_r_46')
// (10, 19, 'sp4_r_v_b_2')
// (10, 19, 'sp4_r_v_b_6')
// (11, 11, 'sp12_h_r_16')
// (11, 11, 'sp4_h_r_0')
// (11, 11, 'sp4_v_t_37')
// (11, 11, 'sp4_v_t_43')
// (11, 12, 'sp4_v_b_37')
// (11, 12, 'sp4_v_b_43')
// (11, 13, 'sp4_v_b_24')
// (11, 13, 'sp4_v_b_30')
// (11, 14, 'sp4_v_b_13')
// (11, 14, 'sp4_v_b_19')
// (11, 15, 'sp4_h_r_19')
// (11, 15, 'sp4_h_r_2')
// (11, 15, 'sp4_v_b_0')
// (11, 15, 'sp4_v_b_6')
// (11, 15, 'sp4_v_t_39')
// (11, 15, 'sp4_v_t_43')
// (11, 16, 'sp4_v_b_39')
// (11, 16, 'sp4_v_b_43')
// (11, 17, 'local_g2_6')
// (11, 17, 'lutff_1/in_1')
// (11, 17, 'sp4_v_b_26')
// (11, 17, 'sp4_v_b_30')
// (11, 18, 'sp4_v_b_15')
// (11, 18, 'sp4_v_b_19')
// (11, 19, 'sp4_h_l_46')
// (11, 19, 'sp4_h_r_15')
// (11, 19, 'sp4_v_b_2')
// (11, 19, 'sp4_v_b_6')
// (12, 11, 'sp12_h_r_19')
// (12, 11, 'sp4_h_r_13')
// (12, 15, 'sp4_h_r_15')
// (12, 15, 'sp4_h_r_30')
// (12, 19, 'sp4_h_r_26')
// (12, 19, 'sp4_h_r_3')
// (13, 11, 'sp12_h_r_20')
// (13, 11, 'sp4_h_r_24')
// (13, 12, 'sp4_r_v_b_36')
// (13, 13, 'sp4_r_v_b_25')
// (13, 14, 'sp4_r_v_b_12')
// (13, 15, 'local_g2_2')
// (13, 15, 'lutff_global/cen')
// (13, 15, 'sp4_h_r_26')
// (13, 15, 'sp4_h_r_43')
// (13, 15, 'sp4_r_v_b_1')
// (13, 16, 'sp4_r_v_b_36')
// (13, 16, 'sp4_r_v_b_44')
// (13, 17, 'local_g0_2')
// (13, 17, 'lutff_4/in_0')
// (13, 17, 'sp4_r_v_b_25')
// (13, 17, 'sp4_r_v_b_33')
// (13, 18, 'sp4_r_v_b_12')
// (13, 18, 'sp4_r_v_b_20')
// (13, 19, 'sp4_h_r_14')
// (13, 19, 'sp4_h_r_39')
// (13, 19, 'sp4_r_v_b_1')
// (13, 19, 'sp4_r_v_b_9')
// (13, 20, 'sp4_r_v_b_41')
// (13, 21, 'local_g1_4')
// (13, 21, 'lutff_7/in_2')
// (13, 21, 'sp4_r_v_b_28')
// (13, 22, 'sp4_r_v_b_17')
// (13, 23, 'sp4_r_v_b_4')
// (14, 1, 'neigh_op_bnr_2')
// (14, 1, 'neigh_op_bnr_6')
// (14, 8, 'sp4_r_v_b_37')
// (14, 9, 'sp4_r_v_b_24')
// (14, 10, 'sp4_r_v_b_13')
// (14, 11, 'sp12_h_r_23')
// (14, 11, 'sp4_h_r_1')
// (14, 11, 'sp4_h_r_37')
// (14, 11, 'sp4_r_v_b_0')
// (14, 11, 'sp4_v_t_36')
// (14, 12, 'local_g2_5')
// (14, 12, 'local_g3_5')
// (14, 12, 'lutff_4/in_2')
// (14, 12, 'lutff_5/in_0')
// (14, 12, 'sp4_r_v_b_37')
// (14, 12, 'sp4_r_v_b_45')
// (14, 12, 'sp4_v_b_36')
// (14, 13, 'sp4_r_v_b_24')
// (14, 13, 'sp4_r_v_b_32')
// (14, 13, 'sp4_v_b_25')
// (14, 14, 'sp4_r_v_b_13')
// (14, 14, 'sp4_r_v_b_21')
// (14, 14, 'sp4_v_b_12')
// (14, 15, 'sp4_h_l_43')
// (14, 15, 'sp4_h_r_39')
// (14, 15, 'sp4_r_v_b_0')
// (14, 15, 'sp4_r_v_b_8')
// (14, 15, 'sp4_v_b_1')
// (14, 15, 'sp4_v_t_36')
// (14, 15, 'sp4_v_t_44')
// (14, 16, 'local_g2_6')
// (14, 16, 'lutff_5/in_1')
// (14, 16, 'lutff_6/in_0')
// (14, 16, 'sp4_r_v_b_38')
// (14, 16, 'sp4_v_b_36')
// (14, 16, 'sp4_v_b_44')
// (14, 17, 'sp4_r_v_b_27')
// (14, 17, 'sp4_v_b_25')
// (14, 17, 'sp4_v_b_33')
// (14, 18, 'sp4_r_v_b_14')
// (14, 18, 'sp4_v_b_12')
// (14, 18, 'sp4_v_b_20')
// (14, 19, 'sp4_h_l_39')
// (14, 19, 'sp4_h_r_27')
// (14, 19, 'sp4_r_v_b_3')
// (14, 19, 'sp4_v_b_1')
// (14, 19, 'sp4_v_b_9')
// (14, 19, 'sp4_v_t_41')
// (14, 20, 'sp4_v_b_41')
// (14, 21, 'sp4_v_b_28')
// (14, 22, 'sp4_v_b_17')
// (14, 23, 'sp4_v_b_4')
// (15, 0, 'io_1/D_IN_0')
// (15, 0, 'io_1/PAD')
// (15, 0, 'span12_vert_12')
// (15, 0, 'span12_vert_20')
// (15, 0, 'span4_horz_r_2')
// (15, 1, 'neigh_op_bot_2')
// (15, 1, 'neigh_op_bot_6')
// (15, 1, 'sp12_v_b_12')
// (15, 1, 'sp12_v_b_20')
// (15, 2, 'sp12_v_b_11')
// (15, 2, 'sp12_v_b_19')
// (15, 3, 'sp12_v_b_16')
// (15, 3, 'sp12_v_b_8')
// (15, 4, 'sp12_v_b_15')
// (15, 4, 'sp12_v_b_7')
// (15, 5, 'sp12_v_b_12')
// (15, 5, 'sp12_v_b_4')
// (15, 6, 'sp12_v_b_11')
// (15, 6, 'sp12_v_b_3')
// (15, 7, 'sp12_v_b_0')
// (15, 7, 'sp12_v_b_8')
// (15, 7, 'sp12_v_t_23')
// (15, 7, 'sp4_v_t_37')
// (15, 8, 'sp12_v_b_23')
// (15, 8, 'sp12_v_b_7')
// (15, 8, 'sp4_v_b_37')
// (15, 9, 'sp12_v_b_20')
// (15, 9, 'sp12_v_b_4')
// (15, 9, 'sp4_v_b_24')
// (15, 10, 'sp12_v_b_19')
// (15, 10, 'sp12_v_b_3')
// (15, 10, 'sp4_v_b_13')
// (15, 11, 'sp12_h_l_23')
// (15, 11, 'sp12_h_r_0')
// (15, 11, 'sp12_v_b_0')
// (15, 11, 'sp12_v_b_16')
// (15, 11, 'sp4_h_l_37')
// (15, 11, 'sp4_h_r_12')
// (15, 11, 'sp4_v_b_0')
// (15, 11, 'sp4_v_t_37')
// (15, 11, 'sp4_v_t_45')
// (15, 12, 'sp12_v_b_15')
// (15, 12, 'sp4_v_b_37')
// (15, 12, 'sp4_v_b_45')
// (15, 13, 'sp12_v_b_12')
// (15, 13, 'sp4_v_b_24')
// (15, 13, 'sp4_v_b_32')
// (15, 14, 'sp12_v_b_11')
// (15, 14, 'sp4_v_b_13')
// (15, 14, 'sp4_v_b_21')
// (15, 15, 'sp12_v_b_8')
// (15, 15, 'sp4_h_l_39')
// (15, 15, 'sp4_h_r_2')
// (15, 15, 'sp4_v_b_0')
// (15, 15, 'sp4_v_b_8')
// (15, 15, 'sp4_v_t_38')
// (15, 16, 'sp12_v_b_7')
// (15, 16, 'sp4_v_b_38')
// (15, 17, 'sp12_v_b_4')
// (15, 17, 'sp4_v_b_27')
// (15, 18, 'sp12_v_b_3')
// (15, 18, 'sp4_v_b_14')
// (15, 19, 'sp12_h_r_0')
// (15, 19, 'sp12_v_b_0')
// (15, 19, 'sp4_h_r_38')
// (15, 19, 'sp4_v_b_3')
// (15, 20, 'sp4_h_r_2')
// (15, 20, 'sp4_r_v_b_45')
// (15, 21, 'sp4_r_v_b_32')
// (15, 22, 'sp4_r_v_b_21')
// (15, 23, 'sp4_r_v_b_8')
// (16, 0, 'span4_horz_r_6')
// (16, 1, 'neigh_op_bnl_2')
// (16, 1, 'neigh_op_bnl_6')
// (16, 11, 'sp12_h_r_3')
// (16, 11, 'sp4_h_r_25')
// (16, 15, 'local_g1_7')
// (16, 15, 'lutff_7/in_1')
// (16, 15, 'sp4_h_r_15')
// (16, 19, 'sp12_h_r_3')
// (16, 19, 'sp4_h_l_38')
// (16, 19, 'sp4_h_r_3')
// (16, 19, 'sp4_v_t_45')
// (16, 20, 'local_g0_7')
// (16, 20, 'lutff_0/in_1')
// (16, 20, 'sp4_h_r_15')
// (16, 20, 'sp4_v_b_45')
// (16, 21, 'sp4_v_b_32')
// (16, 22, 'local_g0_5')
// (16, 22, 'lutff_4/in_1')
// (16, 22, 'lutff_5/in_0')
// (16, 22, 'sp4_v_b_21')
// (16, 23, 'sp4_h_r_2')
// (16, 23, 'sp4_v_b_8')
// (17, 0, 'span4_horz_r_10')
// (17, 11, 'sp12_h_r_4')
// (17, 11, 'sp4_h_r_36')
// (17, 15, 'sp4_h_r_26')
// (17, 19, 'sp12_h_r_4')
// (17, 19, 'sp4_h_r_14')
// (17, 20, 'sp4_h_r_26')
// (17, 23, 'sp4_h_r_15')
// (18, 0, 'span4_horz_r_14')
// (18, 1, 'sp4_r_v_b_37')
// (18, 2, 'sp4_r_v_b_24')
// (18, 3, 'sp4_r_v_b_13')
// (18, 4, 'sp4_r_v_b_0')
// (18, 5, 'sp4_r_v_b_38')
// (18, 6, 'sp4_r_v_b_27')
// (18, 7, 'sp4_r_v_b_14')
// (18, 8, 'sp4_r_v_b_3')
// (18, 9, 'sp4_r_v_b_43')
// (18, 10, 'sp4_r_v_b_30')
// (18, 11, 'sp12_h_r_7')
// (18, 11, 'sp4_h_l_36')
// (18, 11, 'sp4_r_v_b_19')
// (18, 12, 'sp4_r_v_b_6')
// (18, 13, 'sp4_r_v_b_44')
// (18, 14, 'sp4_r_v_b_33')
// (18, 15, 'sp4_h_r_39')
// (18, 15, 'sp4_r_v_b_20')
// (18, 16, 'sp4_r_v_b_9')
// (18, 17, 'sp4_r_v_b_44')
// (18, 18, 'sp4_r_v_b_33')
// (18, 19, 'sp12_h_r_7')
// (18, 19, 'sp4_h_r_27')
// (18, 19, 'sp4_r_v_b_20')
// (18, 20, 'sp4_h_r_39')
// (18, 20, 'sp4_r_v_b_9')
// (18, 21, 'sp4_r_v_b_40')
// (18, 22, 'local_g0_5')
// (18, 22, 'lutff_0/in_1')
// (18, 22, 'lutff_5/in_2')
// (18, 22, 'lutff_6/in_1')
// (18, 22, 'lutff_7/in_2')
// (18, 22, 'sp4_r_v_b_29')
// (18, 23, 'sp4_h_r_26')
// (18, 23, 'sp4_r_v_b_16')
// (18, 24, 'sp4_r_v_b_5')
// (19, 0, 'span4_horz_l_14')
// (19, 0, 'span4_horz_r_2')
// (19, 0, 'span4_vert_37')
// (19, 1, 'sp4_v_b_37')
// (19, 2, 'sp4_v_b_24')
// (19, 3, 'sp4_v_b_13')
// (19, 4, 'sp4_v_b_0')
// (19, 4, 'sp4_v_t_38')
// (19, 5, 'sp4_v_b_38')
// (19, 6, 'sp4_v_b_27')
// (19, 7, 'sp4_v_b_14')
// (19, 8, 'sp4_v_b_3')
// (19, 8, 'sp4_v_t_43')
// (19, 9, 'sp4_v_b_43')
// (19, 10, 'sp4_v_b_30')
// (19, 11, 'sp12_h_r_8')
// (19, 11, 'sp4_v_b_19')
// (19, 12, 'local_g0_6')
// (19, 12, 'lutff_4/in_2')
// (19, 12, 'sp4_v_b_6')
// (19, 12, 'sp4_v_t_44')
// (19, 13, 'sp4_v_b_44')
// (19, 14, 'sp4_v_b_33')
// (19, 15, 'sp4_h_l_39')
// (19, 15, 'sp4_v_b_20')
// (19, 16, 'sp4_v_b_9')
// (19, 16, 'sp4_v_t_44')
// (19, 17, 'sp4_v_b_44')
// (19, 18, 'sp4_v_b_33')
// (19, 19, 'sp12_h_r_8')
// (19, 19, 'sp4_h_r_38')
// (19, 19, 'sp4_v_b_20')
// (19, 20, 'local_g1_1')
// (19, 20, 'lutff_0/in_2')
// (19, 20, 'lutff_1/in_1')
// (19, 20, 'lutff_2/in_2')
// (19, 20, 'lutff_3/in_1')
// (19, 20, 'lutff_4/in_2')
// (19, 20, 'sp4_h_l_39')
// (19, 20, 'sp4_v_b_9')
// (19, 20, 'sp4_v_t_40')
// (19, 21, 'sp4_v_b_40')
// (19, 22, 'sp4_v_b_29')
// (19, 23, 'local_g3_7')
// (19, 23, 'lutff_0/in_2')
// (19, 23, 'lutff_1/in_1')
// (19, 23, 'lutff_2/in_2')
// (19, 23, 'lutff_3/in_1')
// (19, 23, 'lutff_4/in_2')
// (19, 23, 'lutff_5/in_1')
// (19, 23, 'lutff_6/in_2')
// (19, 23, 'lutff_7/in_1')
// (19, 23, 'sp4_h_r_39')
// (19, 23, 'sp4_v_b_16')
// (19, 24, 'sp4_v_b_5')
// (20, 0, 'fabout')
// (20, 0, 'local_g1_6')
// (20, 0, 'span4_horz_r_6')
// (20, 11, 'sp12_h_r_11')
// (20, 19, 'sp12_h_r_11')
// (20, 19, 'sp4_h_l_38')
// (20, 23, 'sp4_h_l_39')
// (21, 0, 'span4_horz_r_10')
// (21, 11, 'sp12_h_r_12')
// (21, 19, 'sp12_h_r_12')
// (22, 0, 'span4_horz_r_14')
// (22, 11, 'sp12_h_r_15')
// (22, 19, 'sp12_h_r_15')
// (23, 0, 'span4_horz_l_14')
// (23, 11, 'sp12_h_r_16')
// (23, 19, 'sp12_h_r_16')
// (24, 11, 'sp12_h_r_19')
// (24, 19, 'sp12_h_r_19')
// (25, 11, 'sp12_h_r_20')
// (25, 19, 'sp12_h_r_20')
// (26, 11, 'sp12_h_r_23')
// (26, 19, 'sp12_h_r_23')
// (27, 11, 'sp12_h_l_23')
// (27, 19, 'sp12_h_l_23')

reg io_0_27_1 = 0;
// (0, 27, 'io_1/D_OUT_0')
// (0, 27, 'io_1/PAD')
// (0, 27, 'local_g0_7')
// (0, 27, 'span12_horz_23')
// (1, 15, 'sp12_h_r_0')
// (1, 15, 'sp12_v_t_23')
// (1, 16, 'sp12_v_b_23')
// (1, 17, 'sp12_v_b_20')
// (1, 18, 'sp12_v_b_19')
// (1, 19, 'sp12_v_b_16')
// (1, 20, 'sp12_v_b_15')
// (1, 21, 'sp12_v_b_12')
// (1, 22, 'sp12_v_b_11')
// (1, 23, 'sp12_v_b_8')
// (1, 24, 'sp12_v_b_7')
// (1, 25, 'sp12_v_b_4')
// (1, 26, 'sp12_v_b_3')
// (1, 27, 'sp12_h_l_23')
// (1, 27, 'sp12_v_b_0')
// (2, 15, 'sp12_h_r_3')
// (3, 15, 'sp12_h_r_4')
// (4, 15, 'sp12_h_r_7')
// (5, 15, 'sp12_h_r_8')
// (6, 13, 'sp4_r_v_b_44')
// (6, 14, 'neigh_op_tnr_2')
// (6, 14, 'sp4_r_v_b_33')
// (6, 15, 'neigh_op_rgt_2')
// (6, 15, 'sp12_h_r_11')
// (6, 15, 'sp4_r_v_b_20')
// (6, 16, 'neigh_op_bnr_2')
// (6, 16, 'sp4_r_v_b_9')
// (7, 12, 'sp4_v_t_44')
// (7, 13, 'sp4_v_b_44')
// (7, 14, 'neigh_op_top_2')
// (7, 14, 'sp4_v_b_33')
// (7, 15, 'lutff_2/out')
// (7, 15, 'sp12_h_r_12')
// (7, 15, 'sp4_v_b_20')
// (7, 16, 'neigh_op_bot_2')
// (7, 16, 'sp4_h_r_9')
// (7, 16, 'sp4_v_b_9')
// (8, 14, 'neigh_op_tnl_2')
// (8, 15, 'neigh_op_lft_2')
// (8, 15, 'sp12_h_r_15')
// (8, 16, 'neigh_op_bnl_2')
// (8, 16, 'sp4_h_r_20')
// (9, 15, 'sp12_h_r_16')
// (9, 16, 'sp4_h_r_33')
// (10, 15, 'sp12_h_r_19')
// (10, 16, 'sp4_h_r_44')
// (11, 15, 'sp12_h_r_20')
// (11, 16, 'local_g0_0')
// (11, 16, 'lutff_0/in_2')
// (11, 16, 'sp4_h_l_44')
// (11, 16, 'sp4_h_r_0')
// (12, 15, 'sp12_h_r_23')
// (12, 16, 'local_g0_5')
// (12, 16, 'lutff_5/in_2')
// (12, 16, 'sp4_h_r_13')
// (13, 15, 'sp12_h_l_23')
// (13, 16, 'sp4_h_r_24')
// (14, 16, 'sp4_h_r_37')
// (15, 16, 'sp4_h_l_37')

wire io_0_30_0;
// (0, 27, 'span4_horz_19')
// (0, 27, 'span4_vert_t_15')
// (0, 28, 'span4_vert_b_15')
// (0, 29, 'span4_vert_b_11')
// (0, 30, 'io_0/D_OUT_0')
// (0, 30, 'io_0/PAD')
// (0, 30, 'local_g1_7')
// (0, 30, 'span4_vert_b_7')
// (0, 31, 'span4_vert_b_3')
// (1, 27, 'sp4_h_r_30')
// (2, 27, 'sp4_h_r_43')
// (2, 28, 'sp4_r_v_b_37')
// (2, 29, 'sp4_r_v_b_24')
// (2, 30, 'sp4_r_v_b_13')
// (2, 31, 'sp4_r_v_b_0')
// (3, 19, 'sp12_h_r_0')
// (3, 19, 'sp12_v_t_23')
// (3, 20, 'sp12_v_b_23')
// (3, 21, 'sp12_v_b_20')
// (3, 22, 'sp12_v_b_19')
// (3, 23, 'sp12_v_b_16')
// (3, 24, 'sp12_v_b_15')
// (3, 25, 'sp12_v_b_12')
// (3, 26, 'sp12_v_b_11')
// (3, 27, 'sp12_v_b_8')
// (3, 27, 'sp4_h_l_43')
// (3, 27, 'sp4_v_t_37')
// (3, 28, 'sp12_v_b_7')
// (3, 28, 'sp4_v_b_37')
// (3, 29, 'sp12_v_b_4')
// (3, 29, 'sp4_v_b_24')
// (3, 30, 'sp12_v_b_3')
// (3, 30, 'sp4_v_b_13')
// (3, 31, 'sp12_v_b_0')
// (3, 31, 'sp4_v_b_0')
// (4, 19, 'sp12_h_r_3')
// (5, 19, 'sp12_h_r_4')
// (6, 19, 'sp12_h_r_7')
// (7, 19, 'sp12_h_r_8')
// (8, 18, 'neigh_op_tnr_2')
// (8, 19, 'neigh_op_rgt_2')
// (8, 19, 'sp12_h_r_11')
// (8, 20, 'neigh_op_bnr_2')
// (9, 18, 'neigh_op_top_2')
// (9, 19, 'lutff_2/out')
// (9, 19, 'sp12_h_r_12')
// (9, 20, 'neigh_op_bot_2')
// (10, 18, 'neigh_op_tnl_2')
// (10, 19, 'neigh_op_lft_2')
// (10, 19, 'sp12_h_r_15')
// (10, 20, 'neigh_op_bnl_2')
// (11, 19, 'sp12_h_r_16')
// (12, 19, 'sp12_h_r_19')
// (13, 19, 'sp12_h_r_20')
// (14, 19, 'sp12_h_r_23')
// (15, 19, 'sp12_h_l_23')

wire io_0_28_1;
// (0, 28, 'io_1/D_IN_0')
// (0, 28, 'io_1/PAD')
// (0, 28, 'span12_horz_12')
// (1, 27, 'neigh_op_tnl_2')
// (1, 27, 'neigh_op_tnl_6')
// (1, 28, 'neigh_op_lft_2')
// (1, 28, 'neigh_op_lft_6')
// (1, 28, 'sp12_h_r_15')
// (1, 29, 'neigh_op_bnl_2')
// (1, 29, 'neigh_op_bnl_6')
// (2, 28, 'sp12_h_r_16')
// (3, 28, 'sp12_h_r_19')
// (4, 28, 'sp12_h_r_20')
// (5, 19, 'sp4_r_v_b_43')
// (5, 20, 'local_g0_6')
// (5, 20, 'lutff_1/in_1')
// (5, 20, 'sp4_r_v_b_30')
// (5, 21, 'sp4_r_v_b_19')
// (5, 22, 'sp4_r_v_b_6')
// (5, 28, 'sp12_h_r_23')
// (6, 16, 'sp12_v_t_23')
// (6, 17, 'sp12_v_b_23')
// (6, 18, 'sp12_v_b_20')
// (6, 18, 'sp4_v_t_43')
// (6, 19, 'sp12_v_b_19')
// (6, 19, 'sp4_v_b_43')
// (6, 20, 'sp12_v_b_16')
// (6, 20, 'sp4_v_b_30')
// (6, 21, 'sp12_v_b_15')
// (6, 21, 'sp4_v_b_19')
// (6, 22, 'sp12_v_b_12')
// (6, 22, 'sp4_v_b_6')
// (6, 23, 'sp12_v_b_11')
// (6, 24, 'sp12_v_b_8')
// (6, 25, 'sp12_v_b_7')
// (6, 26, 'sp12_v_b_4')
// (6, 27, 'sp12_v_b_3')
// (6, 28, 'sp12_h_l_23')
// (6, 28, 'sp12_v_b_0')

wire io_28_0_0;
// (1, 8, 'sp12_h_r_1')
// (2, 8, 'sp12_h_r_2')
// (3, 8, 'sp12_h_r_5')
// (4, 8, 'sp12_h_r_6')
// (5, 7, 'neigh_op_tnr_1')
// (5, 8, 'neigh_op_rgt_1')
// (5, 8, 'sp12_h_r_9')
// (5, 9, 'neigh_op_bnr_1')
// (6, 7, 'neigh_op_top_1')
// (6, 8, 'lutff_1/out')
// (6, 8, 'sp12_h_r_10')
// (6, 9, 'neigh_op_bot_1')
// (7, 7, 'neigh_op_tnl_1')
// (7, 8, 'neigh_op_lft_1')
// (7, 8, 'sp12_h_r_13')
// (7, 9, 'neigh_op_bnl_1')
// (8, 8, 'sp12_h_r_14')
// (9, 8, 'sp12_h_r_17')
// (10, 8, 'sp12_h_r_18')
// (11, 8, 'sp12_h_r_21')
// (12, 8, 'sp12_h_r_22')
// (13, 8, 'sp12_h_l_22')
// (13, 8, 'sp12_h_r_1')
// (14, 8, 'sp12_h_r_2')
// (15, 8, 'sp12_h_r_5')
// (16, 8, 'sp12_h_r_6')
// (17, 8, 'sp12_h_r_9')
// (18, 8, 'sp12_h_r_10')
// (19, 8, 'sp12_h_r_13')
// (20, 8, 'sp12_h_r_14')
// (21, 8, 'sp12_h_r_17')
// (22, 8, 'sp12_h_r_18')
// (23, 8, 'sp12_h_r_21')
// (24, 1, 'sp4_r_v_b_31')
// (24, 2, 'sp4_r_v_b_18')
// (24, 3, 'sp4_r_v_b_7')
// (24, 8, 'sp12_h_r_22')
// (25, 0, 'span12_vert_14')
// (25, 0, 'span4_horz_r_1')
// (25, 0, 'span4_vert_31')
// (25, 1, 'sp12_v_b_14')
// (25, 1, 'sp4_v_b_31')
// (25, 2, 'sp12_v_b_13')
// (25, 2, 'sp4_v_b_18')
// (25, 3, 'sp12_v_b_10')
// (25, 3, 'sp4_v_b_7')
// (25, 4, 'sp12_v_b_9')
// (25, 5, 'sp12_v_b_6')
// (25, 6, 'sp12_v_b_5')
// (25, 7, 'sp12_v_b_2')
// (25, 8, 'sp12_h_l_22')
// (25, 8, 'sp12_v_b_1')
// (26, 0, 'span4_horz_r_5')
// (27, 0, 'span4_horz_r_9')
// (28, 0, 'io_0/D_OUT_0')
// (28, 0, 'io_0/PAD')
// (28, 0, 'local_g1_5')
// (28, 0, 'span4_horz_r_13')
// (29, 0, 'span4_horz_l_13')

wire n26;
// (2, 12, 'sp12_h_r_1')
// (3, 12, 'sp12_h_r_2')
// (4, 12, 'sp12_h_r_5')
// (5, 12, 'sp12_h_r_6')
// (6, 11, 'neigh_op_tnr_1')
// (6, 12, 'neigh_op_rgt_1')
// (6, 12, 'sp12_h_r_9')
// (6, 13, 'neigh_op_bnr_1')
// (7, 10, 'sp4_r_v_b_43')
// (7, 11, 'neigh_op_top_1')
// (7, 11, 'sp4_r_v_b_30')
// (7, 12, 'lutff_1/out')
// (7, 12, 'sp12_h_r_10')
// (7, 12, 'sp4_r_v_b_19')
// (7, 13, 'neigh_op_bot_1')
// (7, 13, 'sp4_r_v_b_6')
// (8, 9, 'sp4_v_t_43')
// (8, 10, 'sp4_v_b_43')
// (8, 11, 'neigh_op_tnl_1')
// (8, 11, 'sp4_v_b_30')
// (8, 12, 'neigh_op_lft_1')
// (8, 12, 'sp12_h_r_13')
// (8, 12, 'sp4_v_b_19')
// (8, 13, 'neigh_op_bnl_1')
// (8, 13, 'sp4_h_r_6')
// (8, 13, 'sp4_v_b_6')
// (9, 12, 'sp12_h_r_14')
// (9, 13, 'local_g1_3')
// (9, 13, 'lutff_global/cen')
// (9, 13, 'sp4_h_r_19')
// (10, 12, 'sp12_h_r_17')
// (10, 13, 'sp4_h_r_30')
// (11, 12, 'local_g0_2')
// (11, 12, 'lutff_global/cen')
// (11, 12, 'sp12_h_r_18')
// (11, 13, 'sp4_h_r_43')
// (12, 12, 'sp12_h_r_21')
// (12, 13, 'sp4_h_l_43')
// (13, 12, 'sp12_h_r_22')
// (14, 12, 'sp12_h_l_22')

reg n27 = 0;
// (2, 17, 'sp12_h_r_1')
// (3, 17, 'sp12_h_r_2')
// (4, 16, 'neigh_op_tnr_7')
// (4, 17, 'neigh_op_rgt_7')
// (4, 17, 'sp12_h_r_5')
// (4, 18, 'neigh_op_bnr_7')
// (5, 16, 'neigh_op_top_7')
// (5, 17, 'local_g3_7')
// (5, 17, 'lutff_7/in_1')
// (5, 17, 'lutff_7/out')
// (5, 17, 'sp12_h_r_6')
// (5, 18, 'neigh_op_bot_7')
// (6, 16, 'neigh_op_tnl_7')
// (6, 17, 'neigh_op_lft_7')
// (6, 17, 'sp12_h_r_9')
// (6, 18, 'neigh_op_bnl_7')
// (7, 17, 'sp12_h_r_10')
// (8, 17, 'sp12_h_r_13')
// (9, 17, 'sp12_h_r_14')
// (10, 17, 'sp12_h_r_17')
// (11, 17, 'sp12_h_r_18')
// (12, 17, 'sp12_h_r_21')
// (12, 17, 'sp4_h_r_10')
// (13, 17, 'sp12_h_r_22')
// (13, 17, 'sp4_h_r_23')
// (14, 17, 'sp12_h_l_22')
// (14, 17, 'sp4_h_r_34')
// (15, 17, 'sp4_h_r_47')
// (15, 18, 'sp4_r_v_b_38')
// (15, 19, 'sp4_r_v_b_27')
// (15, 20, 'sp4_r_v_b_14')
// (15, 21, 'sp4_r_v_b_3')
// (15, 22, 'sp4_r_v_b_38')
// (15, 23, 'sp4_r_v_b_27')
// (15, 24, 'sp4_r_v_b_14')
// (15, 25, 'sp4_r_v_b_3')
// (16, 17, 'sp4_h_l_47')
// (16, 17, 'sp4_v_t_38')
// (16, 18, 'sp4_v_b_38')
// (16, 19, 'sp4_v_b_27')
// (16, 20, 'sp4_v_b_14')
// (16, 21, 'sp4_v_b_3')
// (16, 21, 'sp4_v_t_38')
// (16, 22, 'local_g3_6')
// (16, 22, 'lutff_0/in_1')
// (16, 22, 'sp4_v_b_38')
// (16, 23, 'sp4_v_b_27')
// (16, 24, 'sp4_v_b_14')
// (16, 25, 'sp4_v_b_3')

reg n28 = 0;
// (2, 18, 'sp12_h_r_0')
// (2, 19, 'sp4_h_r_5')
// (3, 18, 'sp12_h_r_3')
// (3, 19, 'sp4_h_r_16')
// (4, 12, 'sp12_h_r_0')
// (4, 18, 'sp12_h_r_4')
// (4, 19, 'sp4_h_r_29')
// (5, 12, 'sp12_h_r_3')
// (5, 16, 'sp4_r_v_b_37')
// (5, 17, 'local_g0_0')
// (5, 17, 'local_g1_0')
// (5, 17, 'lutff_0/in_0')
// (5, 17, 'lutff_1/in_0')
// (5, 17, 'lutff_2/in_0')
// (5, 17, 'lutff_3/in_0')
// (5, 17, 'lutff_4/in_0')
// (5, 17, 'lutff_5/in_0')
// (5, 17, 'lutff_6/in_0')
// (5, 17, 'lutff_7/in_0')
// (5, 17, 'sp4_r_v_b_24')
// (5, 18, 'local_g1_7')
// (5, 18, 'local_g2_5')
// (5, 18, 'lutff_0/in_0')
// (5, 18, 'lutff_1/in_0')
// (5, 18, 'lutff_2/in_0')
// (5, 18, 'lutff_3/in_0')
// (5, 18, 'lutff_4/in_0')
// (5, 18, 'lutff_5/in_0')
// (5, 18, 'lutff_6/in_0')
// (5, 18, 'lutff_7/in_0')
// (5, 18, 'sp12_h_r_7')
// (5, 18, 'sp4_r_v_b_13')
// (5, 19, 'local_g1_0')
// (5, 19, 'local_g2_0')
// (5, 19, 'lutff_0/in_0')
// (5, 19, 'lutff_1/in_0')
// (5, 19, 'lutff_2/in_0')
// (5, 19, 'sp4_h_r_40')
// (5, 19, 'sp4_r_v_b_0')
// (6, 12, 'sp12_h_r_4')
// (6, 15, 'sp4_h_r_0')
// (6, 15, 'sp4_v_t_37')
// (6, 16, 'sp4_v_b_37')
// (6, 17, 'sp4_v_b_24')
// (6, 18, 'sp12_h_r_8')
// (6, 18, 'sp4_v_b_13')
// (6, 19, 'sp4_h_l_40')
// (6, 19, 'sp4_v_b_0')
// (7, 12, 'sp12_h_r_7')
// (7, 15, 'sp4_h_r_13')
// (7, 18, 'sp12_h_r_11')
// (8, 12, 'sp12_h_r_8')
// (8, 15, 'sp4_h_r_24')
// (8, 18, 'sp12_h_r_12')
// (9, 12, 'sp12_h_r_11')
// (9, 15, 'sp4_h_r_37')
// (9, 18, 'sp12_h_r_15')
// (10, 12, 'sp12_h_r_12')
// (10, 15, 'sp4_h_l_37')
// (10, 15, 'sp4_h_r_9')
// (10, 18, 'sp12_h_r_16')
// (11, 12, 'sp12_h_r_15')
// (11, 15, 'sp4_h_r_20')
// (11, 18, 'sp12_h_r_19')
// (12, 12, 'sp12_h_r_16')
// (12, 15, 'sp4_h_r_33')
// (12, 18, 'sp12_h_r_20')
// (12, 24, 'sp4_h_r_7')
// (13, 11, 'neigh_op_tnr_6')
// (13, 12, 'neigh_op_rgt_6')
// (13, 12, 'sp12_h_r_19')
// (13, 12, 'sp4_r_v_b_44')
// (13, 13, 'neigh_op_bnr_6')
// (13, 13, 'sp4_r_v_b_33')
// (13, 14, 'sp4_r_v_b_20')
// (13, 15, 'sp4_h_r_44')
// (13, 15, 'sp4_r_v_b_9')
// (13, 16, 'sp4_r_v_b_40')
// (13, 17, 'sp4_r_v_b_29')
// (13, 18, 'sp12_h_r_23')
// (13, 18, 'sp4_r_v_b_16')
// (13, 19, 'sp4_r_v_b_5')
// (13, 20, 'sp4_r_v_b_40')
// (13, 21, 'sp4_r_v_b_29')
// (13, 22, 'sp4_r_v_b_16')
// (13, 23, 'sp4_r_v_b_5')
// (13, 24, 'sp4_h_r_18')
// (14, 6, 'sp12_v_t_23')
// (14, 7, 'sp12_v_b_23')
// (14, 8, 'sp12_v_b_20')
// (14, 9, 'sp12_v_b_19')
// (14, 10, 'sp12_v_b_16')
// (14, 11, 'neigh_op_top_6')
// (14, 11, 'sp12_v_b_15')
// (14, 11, 'sp4_v_t_44')
// (14, 12, 'local_g2_6')
// (14, 12, 'lutff_6/in_0')
// (14, 12, 'lutff_6/out')
// (14, 12, 'sp12_h_r_20')
// (14, 12, 'sp12_v_b_12')
// (14, 12, 'sp4_v_b_44')
// (14, 13, 'neigh_op_bot_6')
// (14, 13, 'sp12_v_b_11')
// (14, 13, 'sp4_v_b_33')
// (14, 14, 'sp12_v_b_8')
// (14, 14, 'sp4_v_b_20')
// (14, 15, 'sp12_v_b_7')
// (14, 15, 'sp4_h_l_44')
// (14, 15, 'sp4_v_b_9')
// (14, 15, 'sp4_v_t_40')
// (14, 16, 'sp12_v_b_4')
// (14, 16, 'sp4_v_b_40')
// (14, 17, 'sp12_v_b_3')
// (14, 17, 'sp4_v_b_29')
// (14, 18, 'sp12_h_l_23')
// (14, 18, 'sp12_v_b_0')
// (14, 18, 'sp4_v_b_16')
// (14, 19, 'sp4_v_b_5')
// (14, 19, 'sp4_v_t_40')
// (14, 20, 'sp4_v_b_40')
// (14, 21, 'sp4_v_b_29')
// (14, 22, 'sp4_v_b_16')
// (14, 23, 'sp4_h_r_11')
// (14, 23, 'sp4_v_b_5')
// (14, 24, 'sp4_h_r_31')
// (15, 11, 'neigh_op_tnl_6')
// (15, 12, 'neigh_op_lft_6')
// (15, 12, 'sp12_h_r_23')
// (15, 13, 'neigh_op_bnl_6')
// (15, 17, 'sp4_r_v_b_41')
// (15, 18, 'sp4_r_v_b_28')
// (15, 19, 'sp4_r_v_b_17')
// (15, 20, 'sp4_r_v_b_4')
// (15, 21, 'sp4_r_v_b_42')
// (15, 22, 'sp4_r_v_b_31')
// (15, 23, 'sp4_h_r_22')
// (15, 23, 'sp4_r_v_b_18')
// (15, 24, 'local_g1_7')
// (15, 24, 'local_g3_2')
// (15, 24, 'lutff_0/in_0')
// (15, 24, 'lutff_1/in_0')
// (15, 24, 'lutff_2/in_0')
// (15, 24, 'lutff_3/in_0')
// (15, 24, 'lutff_4/in_0')
// (15, 24, 'lutff_5/in_0')
// (15, 24, 'lutff_6/in_0')
// (15, 24, 'lutff_7/in_0')
// (15, 24, 'sp4_h_r_42')
// (15, 24, 'sp4_r_v_b_7')
// (15, 25, 'local_g2_6')
// (15, 25, 'local_g3_2')
// (15, 25, 'lutff_0/in_0')
// (15, 25, 'lutff_1/in_0')
// (15, 25, 'lutff_2/in_0')
// (15, 25, 'lutff_3/in_0')
// (15, 25, 'lutff_4/in_0')
// (15, 25, 'lutff_5/in_0')
// (15, 25, 'lutff_6/in_0')
// (15, 25, 'lutff_7/in_0')
// (15, 25, 'sp4_r_v_b_38')
// (15, 25, 'sp4_r_v_b_42')
// (15, 26, 'local_g0_7')
// (15, 26, 'local_g1_3')
// (15, 26, 'lutff_0/in_0')
// (15, 26, 'lutff_1/in_0')
// (15, 26, 'lutff_2/in_0')
// (15, 26, 'sp4_r_v_b_27')
// (15, 26, 'sp4_r_v_b_31')
// (15, 27, 'sp4_r_v_b_14')
// (15, 27, 'sp4_r_v_b_18')
// (15, 28, 'sp4_r_v_b_3')
// (15, 28, 'sp4_r_v_b_7')
// (16, 12, 'sp12_h_l_23')
// (16, 12, 'sp12_v_t_23')
// (16, 13, 'sp12_v_b_23')
// (16, 14, 'sp12_v_b_20')
// (16, 15, 'sp12_v_b_19')
// (16, 16, 'sp12_v_b_16')
// (16, 16, 'sp4_v_t_41')
// (16, 17, 'sp12_v_b_15')
// (16, 17, 'sp4_v_b_41')
// (16, 18, 'sp12_v_b_12')
// (16, 18, 'sp4_v_b_28')
// (16, 19, 'sp12_v_b_11')
// (16, 19, 'sp4_v_b_17')
// (16, 20, 'sp12_v_b_8')
// (16, 20, 'sp4_v_b_4')
// (16, 20, 'sp4_v_t_42')
// (16, 21, 'sp12_v_b_7')
// (16, 21, 'sp4_v_b_42')
// (16, 22, 'local_g3_4')
// (16, 22, 'lutff_3/in_2')
// (16, 22, 'sp12_v_b_4')
// (16, 22, 'sp4_v_b_31')
// (16, 23, 'sp12_v_b_3')
// (16, 23, 'sp4_h_r_35')
// (16, 23, 'sp4_v_b_18')
// (16, 24, 'sp12_v_b_0')
// (16, 24, 'sp4_h_l_42')
// (16, 24, 'sp4_v_b_7')
// (16, 24, 'sp4_v_t_38')
// (16, 24, 'sp4_v_t_42')
// (16, 25, 'sp4_v_b_38')
// (16, 25, 'sp4_v_b_42')
// (16, 26, 'sp4_v_b_27')
// (16, 26, 'sp4_v_b_31')
// (16, 27, 'sp4_v_b_14')
// (16, 27, 'sp4_v_b_18')
// (16, 28, 'sp4_v_b_3')
// (16, 28, 'sp4_v_b_7')
// (17, 23, 'sp4_h_r_46')
// (17, 24, 'sp4_r_v_b_41')
// (17, 25, 'sp4_r_v_b_28')
// (17, 26, 'sp4_r_v_b_17')
// (17, 27, 'sp4_r_v_b_4')
// (18, 23, 'sp4_h_l_46')
// (18, 23, 'sp4_v_t_41')
// (18, 24, 'sp4_v_b_41')
// (18, 25, 'sp4_v_b_28')
// (18, 26, 'local_g1_1')
// (18, 26, 'lutff_0/in_0')
// (18, 26, 'sp4_v_b_17')
// (18, 27, 'sp4_v_b_4')

reg n29 = 0;
// (2, 18, 'sp12_h_r_1')
// (3, 18, 'sp12_h_r_2')
// (4, 17, 'neigh_op_tnr_7')
// (4, 18, 'neigh_op_rgt_7')
// (4, 18, 'sp12_h_r_5')
// (4, 19, 'neigh_op_bnr_7')
// (5, 17, 'neigh_op_top_7')
// (5, 18, 'local_g3_7')
// (5, 18, 'lutff_7/in_1')
// (5, 18, 'lutff_7/out')
// (5, 18, 'sp12_h_r_6')
// (5, 19, 'neigh_op_bot_7')
// (6, 17, 'neigh_op_tnl_7')
// (6, 18, 'neigh_op_lft_7')
// (6, 18, 'sp12_h_r_9')
// (6, 19, 'neigh_op_bnl_7')
// (7, 18, 'sp12_h_r_10')
// (8, 18, 'sp12_h_r_13')
// (9, 18, 'sp12_h_r_14')
// (10, 18, 'sp12_h_r_17')
// (11, 18, 'sp12_h_r_18')
// (12, 18, 'sp12_h_r_21')
// (13, 18, 'sp12_h_r_22')
// (13, 24, 'sp4_r_v_b_40')
// (13, 25, 'sp4_r_v_b_29')
// (13, 26, 'sp4_r_v_b_16')
// (13, 27, 'sp4_r_v_b_5')
// (14, 18, 'sp12_h_l_22')
// (14, 18, 'sp12_v_t_22')
// (14, 19, 'sp12_v_b_22')
// (14, 20, 'sp12_v_b_21')
// (14, 21, 'sp12_v_b_18')
// (14, 22, 'sp12_v_b_17')
// (14, 23, 'sp12_v_b_14')
// (14, 23, 'sp4_h_r_10')
// (14, 23, 'sp4_v_t_40')
// (14, 24, 'sp12_v_b_13')
// (14, 24, 'sp4_v_b_40')
// (14, 25, 'sp12_v_b_10')
// (14, 25, 'sp4_v_b_29')
// (14, 26, 'sp12_v_b_9')
// (14, 26, 'sp4_v_b_16')
// (14, 27, 'sp12_v_b_6')
// (14, 27, 'sp4_v_b_5')
// (14, 28, 'sp12_v_b_5')
// (14, 29, 'sp12_v_b_2')
// (14, 30, 'sp12_v_b_1')
// (15, 23, 'sp4_h_r_23')
// (16, 23, 'sp4_h_r_34')
// (17, 23, 'sp4_h_r_47')
// (18, 23, 'local_g0_2')
// (18, 23, 'lutff_7/in_1')
// (18, 23, 'sp4_h_l_47')
// (18, 23, 'sp4_h_r_10')
// (19, 23, 'sp4_h_r_23')
// (20, 23, 'sp4_h_r_34')
// (21, 23, 'sp4_h_r_47')
// (22, 23, 'sp4_h_l_47')

reg n30 = 0;
// (2, 19, 'sp4_h_r_1')
// (3, 19, 'sp4_h_r_12')
// (4, 18, 'neigh_op_tnr_2')
// (4, 19, 'neigh_op_rgt_2')
// (4, 19, 'sp4_h_r_25')
// (4, 20, 'neigh_op_bnr_2')
// (5, 18, 'neigh_op_top_2')
// (5, 19, 'local_g3_2')
// (5, 19, 'lutff_2/in_1')
// (5, 19, 'lutff_2/out')
// (5, 19, 'sp4_h_r_36')
// (5, 20, 'neigh_op_bot_2')
// (6, 18, 'neigh_op_tnl_2')
// (6, 19, 'neigh_op_lft_2')
// (6, 19, 'sp4_h_l_36')
// (6, 19, 'sp4_h_r_4')
// (6, 20, 'neigh_op_bnl_2')
// (7, 19, 'sp4_h_r_17')
// (8, 19, 'sp4_h_r_28')
// (9, 19, 'sp4_h_r_41')
// (10, 19, 'sp4_h_l_41')
// (10, 19, 'sp4_h_r_0')
// (11, 19, 'sp4_h_r_13')
// (12, 19, 'sp4_h_r_24')
// (13, 19, 'sp4_h_r_37')
// (14, 19, 'sp4_h_l_37')
// (14, 19, 'sp4_h_r_8')
// (15, 19, 'sp4_h_r_21')
// (16, 19, 'sp4_h_r_32')
// (17, 19, 'sp4_h_r_45')
// (17, 20, 'sp4_r_v_b_45')
// (17, 21, 'sp4_r_v_b_32')
// (17, 22, 'sp4_r_v_b_21')
// (17, 23, 'sp4_r_v_b_8')
// (18, 19, 'sp4_h_l_45')
// (18, 19, 'sp4_v_t_45')
// (18, 20, 'sp4_v_b_45')
// (18, 21, 'local_g2_0')
// (18, 21, 'lutff_2/in_2')
// (18, 21, 'sp4_v_b_32')
// (18, 22, 'sp4_v_b_21')
// (18, 23, 'sp4_v_b_8')

reg n31 = 0;
// (2, 21, 'sp12_h_r_0')
// (3, 21, 'sp12_h_r_3')
// (4, 21, 'sp12_h_r_4')
// (5, 21, 'sp12_h_r_7')
// (6, 21, 'sp12_h_r_8')
// (7, 21, 'sp12_h_r_11')
// (8, 21, 'sp12_h_r_12')
// (9, 21, 'sp12_h_r_15')
// (10, 21, 'sp12_h_r_16')
// (11, 21, 'sp12_h_r_19')
// (12, 21, 'local_g1_4')
// (12, 21, 'lutff_4/in_3')
// (12, 21, 'sp12_h_r_20')
// (13, 21, 'sp12_h_r_23')
// (13, 22, 'neigh_op_tnr_2')
// (13, 23, 'neigh_op_rgt_2')
// (13, 24, 'neigh_op_bnr_2')
// (14, 21, 'sp12_h_l_23')
// (14, 21, 'sp12_v_t_23')
// (14, 22, 'neigh_op_top_2')
// (14, 22, 'sp12_v_b_23')
// (14, 23, 'lutff_2/out')
// (14, 23, 'sp12_v_b_20')
// (14, 24, 'neigh_op_bot_2')
// (14, 24, 'sp12_v_b_19')
// (14, 25, 'sp12_v_b_16')
// (14, 26, 'sp12_v_b_15')
// (14, 27, 'sp12_v_b_12')
// (14, 28, 'sp12_v_b_11')
// (14, 29, 'sp12_v_b_8')
// (14, 30, 'sp12_v_b_7')
// (14, 31, 'sp12_v_b_4')
// (14, 32, 'sp12_v_b_3')
// (14, 33, 'span12_vert_0')
// (15, 22, 'neigh_op_tnl_2')
// (15, 23, 'neigh_op_lft_2')
// (15, 24, 'neigh_op_bnl_2')

wire n32;
// (2, 23, 'sp12_h_r_1')
// (3, 23, 'sp12_h_r_2')
// (4, 23, 'sp12_h_r_5')
// (5, 23, 'sp12_h_r_6')
// (6, 23, 'sp12_h_r_9')
// (7, 23, 'sp12_h_r_10')
// (8, 23, 'sp12_h_r_13')
// (9, 14, 'sp12_h_r_1')
// (9, 23, 'sp12_h_r_14')
// (10, 10, 'local_g0_2')
// (10, 10, 'local_g1_2')
// (10, 10, 'lutff_5/in_1')
// (10, 10, 'lutff_6/in_1')
// (10, 10, 'lutff_7/in_1')
// (10, 10, 'sp4_h_r_2')
// (10, 14, 'sp12_h_r_2')
// (10, 15, 'sp4_h_r_0')
// (10, 15, 'sp4_r_v_b_39')
// (10, 16, 'sp4_r_v_b_26')
// (10, 17, 'local_g2_7')
// (10, 17, 'lutff_6/in_1')
// (10, 17, 'lutff_7/in_2')
// (10, 17, 'sp4_r_v_b_15')
// (10, 18, 'sp4_r_v_b_2')
// (10, 23, 'sp12_h_r_17')
// (11, 10, 'sp4_h_r_15')
// (11, 14, 'local_g1_2')
// (11, 14, 'local_g1_5')
// (11, 14, 'lutff_1/in_1')
// (11, 14, 'lutff_2/in_1')
// (11, 14, 'lutff_3/in_1')
// (11, 14, 'lutff_4/in_1')
// (11, 14, 'lutff_5/in_1')
// (11, 14, 'lutff_6/in_1')
// (11, 14, 'lutff_7/in_1')
// (11, 14, 'sp12_h_r_5')
// (11, 14, 'sp4_h_r_2')
// (11, 14, 'sp4_v_t_39')
// (11, 15, 'local_g0_5')
// (11, 15, 'local_g3_7')
// (11, 15, 'lutff_0/in_1')
// (11, 15, 'lutff_1/in_1')
// (11, 15, 'lutff_2/in_1')
// (11, 15, 'lutff_3/in_1')
// (11, 15, 'lutff_4/in_1')
// (11, 15, 'lutff_5/in_1')
// (11, 15, 'lutff_6/in_1')
// (11, 15, 'sp4_h_r_13')
// (11, 15, 'sp4_v_b_39')
// (11, 16, 'sp4_v_b_26')
// (11, 17, 'sp4_v_b_15')
// (11, 18, 'sp4_v_b_2')
// (11, 22, 'sp4_h_r_10')
// (11, 23, 'sp12_h_r_18')
// (12, 10, 'sp4_h_r_26')
// (12, 14, 'sp12_h_r_6')
// (12, 14, 'sp4_h_r_15')
// (12, 15, 'sp4_h_r_24')
// (12, 22, 'local_g0_7')
// (12, 22, 'lutff_0/in_1')
// (12, 22, 'lutff_1/in_2')
// (12, 22, 'lutff_2/in_1')
// (12, 22, 'lutff_3/in_2')
// (12, 22, 'lutff_4/in_1')
// (12, 22, 'lutff_5/in_2')
// (12, 22, 'lutff_6/in_1')
// (12, 22, 'lutff_7/in_2')
// (12, 22, 'sp4_h_r_23')
// (12, 23, 'local_g0_5')
// (12, 23, 'lutff_0/in_1')
// (12, 23, 'lutff_1/in_2')
// (12, 23, 'lutff_2/in_1')
// (12, 23, 'lutff_3/in_2')
// (12, 23, 'lutff_4/in_1')
// (12, 23, 'lutff_5/in_2')
// (12, 23, 'lutff_6/in_1')
// (12, 23, 'lutff_7/in_2')
// (12, 23, 'sp12_h_r_21')
// (13, 10, 'sp4_h_r_39')
// (13, 11, 'sp4_r_v_b_39')
// (13, 12, 'sp4_r_v_b_26')
// (13, 12, 'sp4_r_v_b_42')
// (13, 13, 'neigh_op_tnr_1')
// (13, 13, 'sp4_r_v_b_15')
// (13, 13, 'sp4_r_v_b_31')
// (13, 14, 'neigh_op_rgt_1')
// (13, 14, 'sp12_h_r_9')
// (13, 14, 'sp4_h_r_26')
// (13, 14, 'sp4_r_v_b_18')
// (13, 14, 'sp4_r_v_b_2')
// (13, 15, 'neigh_op_bnr_1')
// (13, 15, 'sp4_h_r_37')
// (13, 15, 'sp4_r_v_b_7')
// (13, 19, 'sp4_r_v_b_38')
// (13, 20, 'sp4_r_v_b_27')
// (13, 21, 'sp4_r_v_b_14')
// (13, 21, 'sp4_r_v_b_36')
// (13, 22, 'sp4_h_r_34')
// (13, 22, 'sp4_r_v_b_25')
// (13, 22, 'sp4_r_v_b_3')
// (13, 23, 'local_g1_6')
// (13, 23, 'lutff_0/in_1')
// (13, 23, 'lutff_1/in_2')
// (13, 23, 'lutff_2/in_1')
// (13, 23, 'lutff_3/in_2')
// (13, 23, 'lutff_4/in_1')
// (13, 23, 'lutff_5/in_2')
// (13, 23, 'lutff_6/in_1')
// (13, 23, 'lutff_7/in_2')
// (13, 23, 'sp12_h_r_22')
// (13, 23, 'sp4_r_v_b_12')
// (13, 23, 'sp4_r_v_b_46')
// (13, 24, 'local_g2_3')
// (13, 24, 'lutff_0/in_1')
// (13, 24, 'lutff_1/in_2')
// (13, 24, 'lutff_2/in_1')
// (13, 24, 'lutff_3/in_2')
// (13, 24, 'lutff_4/in_1')
// (13, 24, 'lutff_5/in_2')
// (13, 24, 'lutff_6/in_1')
// (13, 24, 'lutff_7/in_2')
// (13, 24, 'sp4_r_v_b_1')
// (13, 24, 'sp4_r_v_b_35')
// (13, 25, 'sp4_r_v_b_22')
// (13, 26, 'sp4_r_v_b_11')
// (14, 10, 'sp4_h_l_39')
// (14, 10, 'sp4_h_r_2')
// (14, 10, 'sp4_v_t_39')
// (14, 11, 'sp12_v_t_22')
// (14, 11, 'sp4_v_b_39')
// (14, 11, 'sp4_v_t_42')
// (14, 12, 'sp12_v_b_22')
// (14, 12, 'sp4_v_b_26')
// (14, 12, 'sp4_v_b_42')
// (14, 13, 'neigh_op_top_1')
// (14, 13, 'sp12_v_b_21')
// (14, 13, 'sp4_v_b_15')
// (14, 13, 'sp4_v_b_31')
// (14, 14, 'lutff_1/out')
// (14, 14, 'sp12_h_r_10')
// (14, 14, 'sp12_v_b_18')
// (14, 14, 'sp4_h_r_39')
// (14, 14, 'sp4_v_b_18')
// (14, 14, 'sp4_v_b_2')
// (14, 15, 'neigh_op_bot_1')
// (14, 15, 'sp12_v_b_17')
// (14, 15, 'sp4_h_l_37')
// (14, 15, 'sp4_r_v_b_42')
// (14, 15, 'sp4_v_b_7')
// (14, 16, 'sp12_v_b_14')
// (14, 16, 'sp4_r_v_b_31')
// (14, 17, 'sp12_v_b_13')
// (14, 17, 'sp4_r_v_b_18')
// (14, 18, 'sp12_v_b_10')
// (14, 18, 'sp4_r_v_b_7')
// (14, 18, 'sp4_v_t_38')
// (14, 19, 'sp12_v_b_9')
// (14, 19, 'sp4_r_v_b_47')
// (14, 19, 'sp4_v_b_38')
// (14, 20, 'sp12_v_b_6')
// (14, 20, 'sp4_r_v_b_34')
// (14, 20, 'sp4_v_b_27')
// (14, 20, 'sp4_v_t_36')
// (14, 21, 'sp12_v_b_5')
// (14, 21, 'sp4_r_v_b_23')
// (14, 21, 'sp4_v_b_14')
// (14, 21, 'sp4_v_b_36')
// (14, 22, 'sp12_v_b_2')
// (14, 22, 'sp4_h_r_47')
// (14, 22, 'sp4_r_v_b_10')
// (14, 22, 'sp4_v_b_25')
// (14, 22, 'sp4_v_b_3')
// (14, 22, 'sp4_v_t_46')
// (14, 23, 'sp12_h_l_22')
// (14, 23, 'sp12_v_b_1')
// (14, 23, 'sp4_v_b_12')
// (14, 23, 'sp4_v_b_46')
// (14, 24, 'sp4_h_r_1')
// (14, 24, 'sp4_v_b_1')
// (14, 24, 'sp4_v_b_35')
// (14, 25, 'sp4_v_b_22')
// (14, 26, 'sp4_v_b_11')
// (15, 10, 'sp4_h_r_15')
// (15, 13, 'neigh_op_tnl_1')
// (15, 14, 'neigh_op_lft_1')
// (15, 14, 'sp12_h_r_13')
// (15, 14, 'sp4_h_l_39')
// (15, 14, 'sp4_v_t_42')
// (15, 15, 'neigh_op_bnl_1')
// (15, 15, 'sp4_v_b_42')
// (15, 16, 'sp4_v_b_31')
// (15, 17, 'sp4_v_b_18')
// (15, 18, 'sp4_v_b_7')
// (15, 18, 'sp4_v_t_47')
// (15, 19, 'sp4_v_b_47')
// (15, 20, 'sp4_v_b_34')
// (15, 21, 'sp4_v_b_23')
// (15, 22, 'local_g0_2')
// (15, 22, 'local_g1_2')
// (15, 22, 'lutff_0/in_2')
// (15, 22, 'lutff_1/in_2')
// (15, 22, 'lutff_2/in_2')
// (15, 22, 'lutff_3/in_2')
// (15, 22, 'lutff_4/in_2')
// (15, 22, 'lutff_5/in_1')
// (15, 22, 'lutff_6/in_2')
// (15, 22, 'lutff_7/in_1')
// (15, 22, 'sp4_h_l_47')
// (15, 22, 'sp4_v_b_10')
// (15, 24, 'sp4_h_r_12')
// (16, 10, 'sp4_h_r_26')
// (16, 14, 'sp12_h_r_14')
// (16, 24, 'local_g2_1')
// (16, 24, 'lutff_6/in_3')
// (16, 24, 'sp4_h_r_25')
// (17, 10, 'local_g3_7')
// (17, 10, 'lutff_4/in_0')
// (17, 10, 'lutff_5/in_3')
// (17, 10, 'sp4_h_r_39')
// (17, 14, 'sp12_h_r_17')
// (17, 24, 'local_g2_4')
// (17, 24, 'local_g3_4')
// (17, 24, 'lutff_0/in_2')
// (17, 24, 'lutff_1/in_2')
// (17, 24, 'lutff_2/in_2')
// (17, 24, 'lutff_3/in_1')
// (17, 24, 'lutff_4/in_2')
// (17, 24, 'lutff_5/in_2')
// (17, 24, 'lutff_6/in_2')
// (17, 24, 'lutff_7/in_2')
// (17, 24, 'sp4_h_r_36')
// (18, 10, 'sp4_h_l_39')
// (18, 14, 'sp12_h_r_18')
// (18, 24, 'sp4_h_l_36')
// (19, 14, 'sp12_h_r_21')
// (20, 14, 'sp12_h_r_22')
// (21, 14, 'sp12_h_l_22')

wire io_3_33_1;
// (2, 32, 'neigh_op_tnr_2')
// (2, 32, 'neigh_op_tnr_6')
// (3, 23, 'sp12_h_r_0')
// (3, 23, 'sp12_v_t_23')
// (3, 24, 'sp12_v_b_23')
// (3, 25, 'sp12_v_b_20')
// (3, 26, 'sp12_v_b_19')
// (3, 27, 'sp12_v_b_16')
// (3, 28, 'sp12_v_b_15')
// (3, 29, 'sp12_v_b_12')
// (3, 30, 'sp12_v_b_11')
// (3, 31, 'sp12_v_b_8')
// (3, 32, 'neigh_op_top_2')
// (3, 32, 'neigh_op_top_6')
// (3, 32, 'sp12_v_b_7')
// (3, 33, 'io_1/D_IN_0')
// (3, 33, 'io_1/PAD')
// (3, 33, 'span12_vert_4')
// (4, 23, 'sp12_h_r_3')
// (4, 32, 'neigh_op_tnl_2')
// (4, 32, 'neigh_op_tnl_6')
// (5, 23, 'sp12_h_r_4')
// (6, 23, 'sp12_h_r_7')
// (7, 23, 'sp12_h_r_8')
// (8, 23, 'sp12_h_r_11')
// (9, 23, 'sp12_h_r_12')
// (10, 23, 'sp12_h_r_15')
// (10, 23, 'sp4_h_r_9')
// (11, 23, 'sp12_h_r_16')
// (11, 23, 'sp4_h_r_20')
// (12, 23, 'sp12_h_r_19')
// (12, 23, 'sp4_h_r_33')
// (13, 23, 'sp12_h_r_20')
// (13, 23, 'sp4_h_r_44')
// (14, 23, 'sp12_h_r_23')
// (14, 23, 'sp4_h_l_44')
// (14, 23, 'sp4_h_r_0')
// (15, 23, 'sp12_h_l_23')
// (15, 23, 'sp4_h_r_13')
// (16, 23, 'local_g3_0')
// (16, 23, 'lutff_2/in_3')
// (16, 23, 'sp4_h_r_24')
// (17, 23, 'sp4_h_r_37')
// (18, 23, 'sp4_h_l_37')

reg io_4_0_1 = 0;
// (3, 1, 'sp4_r_v_b_37')
// (3, 2, 'sp4_r_v_b_24')
// (3, 3, 'sp4_r_v_b_13')
// (3, 4, 'sp4_r_v_b_0')
// (3, 5, 'sp4_r_v_b_37')
// (3, 6, 'sp4_r_v_b_24')
// (3, 7, 'sp4_r_v_b_13')
// (3, 8, 'sp4_r_v_b_0')
// (4, 0, 'io_1/D_OUT_0')
// (4, 0, 'io_1/PAD')
// (4, 0, 'local_g0_5')
// (4, 0, 'span4_vert_37')
// (4, 1, 'sp4_v_b_37')
// (4, 2, 'sp4_v_b_24')
// (4, 3, 'sp4_v_b_13')
// (4, 4, 'sp4_v_b_0')
// (4, 4, 'sp4_v_t_37')
// (4, 5, 'sp4_v_b_37')
// (4, 6, 'sp4_v_b_24')
// (4, 7, 'sp4_v_b_13')
// (4, 8, 'sp4_h_r_7')
// (4, 8, 'sp4_v_b_0')
// (5, 8, 'sp4_h_r_18')
// (6, 7, 'neigh_op_tnr_5')
// (6, 8, 'neigh_op_rgt_5')
// (6, 8, 'sp4_h_r_31')
// (6, 9, 'neigh_op_bnr_5')
// (7, 7, 'neigh_op_top_5')
// (7, 8, 'lutff_5/out')
// (7, 8, 'sp4_h_r_42')
// (7, 9, 'neigh_op_bot_5')
// (8, 7, 'neigh_op_tnl_5')
// (8, 8, 'neigh_op_lft_5')
// (8, 8, 'sp4_h_l_42')
// (8, 9, 'neigh_op_bnl_5')

reg n35 = 0;
// (3, 12, 'sp12_h_r_0')
// (4, 12, 'sp12_h_r_3')
// (5, 12, 'sp12_h_r_4')
// (6, 12, 'sp12_h_r_7')
// (7, 12, 'sp12_h_r_8')
// (7, 15, 'sp4_h_r_5')
// (7, 18, 'sp4_h_r_8')
// (8, 12, 'sp12_h_r_11')
// (8, 15, 'sp4_h_r_16')
// (8, 18, 'sp4_h_r_21')
// (9, 12, 'sp12_h_r_12')
// (9, 15, 'local_g3_5')
// (9, 15, 'lutff_6/in_0')
// (9, 15, 'sp4_h_r_29')
// (9, 18, 'local_g3_0')
// (9, 18, 'lutff_0/in_3')
// (9, 18, 'sp4_h_r_32')
// (10, 11, 'neigh_op_tnr_4')
// (10, 11, 'sp4_r_v_b_37')
// (10, 12, 'neigh_op_rgt_4')
// (10, 12, 'sp12_h_r_15')
// (10, 12, 'sp4_r_v_b_24')
// (10, 12, 'sp4_r_v_b_40')
// (10, 13, 'neigh_op_bnr_4')
// (10, 13, 'sp4_r_v_b_13')
// (10, 13, 'sp4_r_v_b_29')
// (10, 14, 'sp4_r_v_b_0')
// (10, 14, 'sp4_r_v_b_16')
// (10, 15, 'sp4_h_r_40')
// (10, 15, 'sp4_r_v_b_45')
// (10, 15, 'sp4_r_v_b_5')
// (10, 16, 'sp4_r_v_b_32')
// (10, 16, 'sp4_r_v_b_45')
// (10, 17, 'sp4_r_v_b_21')
// (10, 17, 'sp4_r_v_b_32')
// (10, 18, 'sp4_h_r_45')
// (10, 18, 'sp4_r_v_b_21')
// (10, 18, 'sp4_r_v_b_8')
// (10, 19, 'local_g2_0')
// (10, 19, 'lutff_4/in_0')
// (10, 19, 'sp4_r_v_b_45')
// (10, 19, 'sp4_r_v_b_8')
// (10, 20, 'local_g0_3')
// (10, 20, 'lutff_2/in_3')
// (10, 20, 'sp4_r_v_b_32')
// (10, 21, 'sp4_r_v_b_21')
// (10, 22, 'sp4_r_v_b_8')
// (11, 10, 'sp4_v_t_37')
// (11, 11, 'neigh_op_top_4')
// (11, 11, 'sp4_v_b_37')
// (11, 11, 'sp4_v_t_40')
// (11, 12, 'lutff_4/out')
// (11, 12, 'sp12_h_r_16')
// (11, 12, 'sp4_h_r_8')
// (11, 12, 'sp4_r_v_b_41')
// (11, 12, 'sp4_v_b_24')
// (11, 12, 'sp4_v_b_40')
// (11, 13, 'local_g1_4')
// (11, 13, 'lutff_2/in_3')
// (11, 13, 'neigh_op_bot_4')
// (11, 13, 'sp4_r_v_b_28')
// (11, 13, 'sp4_v_b_13')
// (11, 13, 'sp4_v_b_29')
// (11, 14, 'sp4_r_v_b_17')
// (11, 14, 'sp4_v_b_0')
// (11, 14, 'sp4_v_b_16')
// (11, 14, 'sp4_v_t_45')
// (11, 15, 'sp4_h_l_40')
// (11, 15, 'sp4_r_v_b_4')
// (11, 15, 'sp4_v_b_45')
// (11, 15, 'sp4_v_b_5')
// (11, 15, 'sp4_v_t_45')
// (11, 16, 'sp4_h_r_6')
// (11, 16, 'sp4_v_b_32')
// (11, 16, 'sp4_v_b_45')
// (11, 17, 'sp4_v_b_21')
// (11, 17, 'sp4_v_b_32')
// (11, 18, 'sp4_h_l_45')
// (11, 18, 'sp4_v_b_21')
// (11, 18, 'sp4_v_b_8')
// (11, 18, 'sp4_v_t_45')
// (11, 19, 'sp4_h_r_2')
// (11, 19, 'sp4_v_b_45')
// (11, 19, 'sp4_v_b_8')
// (11, 20, 'sp4_v_b_32')
// (11, 21, 'sp4_v_b_21')
// (11, 22, 'local_g1_0')
// (11, 22, 'lutff_4/in_3')
// (11, 22, 'sp4_v_b_8')
// (12, 11, 'neigh_op_tnl_4')
// (12, 11, 'sp4_v_t_41')
// (12, 12, 'neigh_op_lft_4')
// (12, 12, 'sp12_h_r_19')
// (12, 12, 'sp4_h_r_21')
// (12, 12, 'sp4_v_b_41')
// (12, 13, 'local_g3_4')
// (12, 13, 'lutff_4/in_3')
// (12, 13, 'neigh_op_bnl_4')
// (12, 13, 'sp4_v_b_28')
// (12, 14, 'sp4_v_b_17')
// (12, 15, 'sp4_h_r_4')
// (12, 15, 'sp4_v_b_4')
// (12, 16, 'sp4_h_r_19')
// (12, 19, 'local_g0_7')
// (12, 19, 'lutff_4/in_3')
// (12, 19, 'sp4_h_r_15')
// (12, 19, 'sp4_h_r_9')
// (13, 12, 'sp12_h_r_20')
// (13, 12, 'sp4_h_r_32')
// (13, 15, 'sp4_h_r_17')
// (13, 16, 'local_g3_6')
// (13, 16, 'lutff_2/in_3')
// (13, 16, 'sp4_h_r_30')
// (13, 19, 'sp4_h_r_20')
// (13, 19, 'sp4_h_r_26')
// (14, 12, 'sp12_h_r_23')
// (14, 12, 'sp4_h_r_45')
// (14, 13, 'local_g2_4')
// (14, 13, 'lutff_4/in_0')
// (14, 13, 'sp4_r_v_b_36')
// (14, 14, 'sp4_r_v_b_25')
// (14, 15, 'sp4_h_r_28')
// (14, 15, 'sp4_r_v_b_12')
// (14, 16, 'sp4_h_r_43')
// (14, 16, 'sp4_r_v_b_1')
// (14, 17, 'sp4_r_v_b_36')
// (14, 18, 'sp4_r_v_b_25')
// (14, 19, 'sp4_h_r_33')
// (14, 19, 'sp4_h_r_39')
// (14, 19, 'sp4_r_v_b_12')
// (14, 20, 'sp4_r_v_b_1')
// (14, 21, 'sp4_r_v_b_41')
// (14, 22, 'sp4_r_v_b_28')
// (14, 23, 'local_g3_1')
// (14, 23, 'lutff_2/in_0')
// (14, 23, 'sp4_r_v_b_17')
// (14, 24, 'sp4_r_v_b_4')
// (15, 12, 'sp12_h_l_23')
// (15, 12, 'sp12_h_r_0')
// (15, 12, 'sp4_h_l_45')
// (15, 12, 'sp4_h_r_8')
// (15, 12, 'sp4_v_t_36')
// (15, 13, 'local_g3_4')
// (15, 13, 'lutff_6/in_1')
// (15, 13, 'sp4_v_b_36')
// (15, 14, 'sp4_v_b_25')
// (15, 15, 'local_g1_4')
// (15, 15, 'lutff_4/in_3')
// (15, 15, 'sp4_h_r_41')
// (15, 15, 'sp4_v_b_12')
// (15, 16, 'sp4_h_l_43')
// (15, 16, 'sp4_h_r_7')
// (15, 16, 'sp4_r_v_b_41')
// (15, 16, 'sp4_v_b_1')
// (15, 16, 'sp4_v_t_36')
// (15, 17, 'local_g3_4')
// (15, 17, 'lutff_4/in_3')
// (15, 17, 'sp4_r_v_b_28')
// (15, 17, 'sp4_v_b_36')
// (15, 18, 'local_g2_1')
// (15, 18, 'lutff_4/in_3')
// (15, 18, 'sp4_r_v_b_17')
// (15, 18, 'sp4_v_b_25')
// (15, 19, 'local_g1_4')
// (15, 19, 'lutff_4/in_3')
// (15, 19, 'sp4_h_l_39')
// (15, 19, 'sp4_h_r_44')
// (15, 19, 'sp4_r_v_b_4')
// (15, 19, 'sp4_v_b_12')
// (15, 20, 'sp4_r_v_b_39')
// (15, 20, 'sp4_v_b_1')
// (15, 20, 'sp4_v_t_41')
// (15, 21, 'sp4_r_v_b_26')
// (15, 21, 'sp4_v_b_41')
// (15, 22, 'sp4_r_v_b_15')
// (15, 22, 'sp4_v_b_28')
// (15, 23, 'sp4_r_v_b_2')
// (15, 23, 'sp4_v_b_17')
// (15, 24, 'sp4_v_b_4')
// (16, 12, 'sp12_h_r_3')
// (16, 12, 'sp4_h_r_21')
// (16, 12, 'sp4_h_r_3')
// (16, 15, 'sp4_h_l_41')
// (16, 15, 'sp4_v_t_41')
// (16, 16, 'local_g1_2')
// (16, 16, 'lutff_4/in_3')
// (16, 16, 'sp4_h_r_18')
// (16, 16, 'sp4_v_b_41')
// (16, 17, 'local_g3_4')
// (16, 17, 'lutff_4/in_3')
// (16, 17, 'sp4_v_b_28')
// (16, 18, 'local_g0_1')
// (16, 18, 'lutff_4/in_1')
// (16, 18, 'sp4_v_b_17')
// (16, 19, 'local_g1_4')
// (16, 19, 'lutff_2/in_3')
// (16, 19, 'sp4_h_l_44')
// (16, 19, 'sp4_v_b_4')
// (16, 19, 'sp4_v_t_39')
// (16, 20, 'sp4_v_b_39')
// (16, 21, 'local_g3_2')
// (16, 21, 'lutff_2/in_3')
// (16, 21, 'sp4_v_b_26')
// (16, 22, 'sp4_v_b_15')
// (16, 23, 'sp4_v_b_2')
// (17, 12, 'sp12_h_r_4')
// (17, 12, 'sp4_h_r_14')
// (17, 12, 'sp4_h_r_32')
// (17, 16, 'sp4_h_r_31')
// (18, 9, 'sp4_r_v_b_39')
// (18, 10, 'sp4_r_v_b_26')
// (18, 11, 'sp4_r_v_b_15')
// (18, 12, 'local_g2_5')
// (18, 12, 'lutff_4/in_3')
// (18, 12, 'sp12_h_r_7')
// (18, 12, 'sp4_h_r_27')
// (18, 12, 'sp4_h_r_45')
// (18, 12, 'sp4_h_r_5')
// (18, 12, 'sp4_r_v_b_2')
// (18, 13, 'sp4_r_v_b_45')
// (18, 14, 'sp4_r_v_b_32')
// (18, 15, 'sp4_r_v_b_21')
// (18, 16, 'sp4_h_r_42')
// (18, 16, 'sp4_r_v_b_8')
// (18, 17, 'sp4_r_v_b_41')
// (18, 17, 'sp4_r_v_b_45')
// (18, 18, 'sp4_r_v_b_28')
// (18, 18, 'sp4_r_v_b_32')
// (18, 19, 'sp4_r_v_b_17')
// (18, 19, 'sp4_r_v_b_21')
// (18, 20, 'local_g2_0')
// (18, 20, 'lutff_6/in_0')
// (18, 20, 'sp4_r_v_b_4')
// (18, 20, 'sp4_r_v_b_8')
// (19, 8, 'sp4_v_t_39')
// (19, 9, 'sp4_r_v_b_44')
// (19, 9, 'sp4_v_b_39')
// (19, 10, 'local_g3_2')
// (19, 10, 'lutff_4/in_3')
// (19, 10, 'sp4_r_v_b_33')
// (19, 10, 'sp4_v_b_26')
// (19, 11, 'local_g0_7')
// (19, 11, 'lutff_4/in_3')
// (19, 11, 'sp4_r_v_b_20')
// (19, 11, 'sp4_v_b_15')
// (19, 12, 'sp12_h_r_8')
// (19, 12, 'sp4_h_l_45')
// (19, 12, 'sp4_h_r_16')
// (19, 12, 'sp4_h_r_38')
// (19, 12, 'sp4_r_v_b_9')
// (19, 12, 'sp4_v_b_2')
// (19, 12, 'sp4_v_t_45')
// (19, 13, 'sp4_r_v_b_45')
// (19, 13, 'sp4_v_b_45')
// (19, 14, 'sp4_r_v_b_32')
// (19, 14, 'sp4_v_b_32')
// (19, 15, 'sp4_r_v_b_21')
// (19, 15, 'sp4_v_b_21')
// (19, 16, 'local_g1_0')
// (19, 16, 'lutff_4/in_3')
// (19, 16, 'sp4_h_l_42')
// (19, 16, 'sp4_r_v_b_8')
// (19, 16, 'sp4_v_b_8')
// (19, 16, 'sp4_v_t_41')
// (19, 16, 'sp4_v_t_45')
// (19, 17, 'sp4_r_v_b_45')
// (19, 17, 'sp4_v_b_41')
// (19, 17, 'sp4_v_b_45')
// (19, 18, 'local_g3_4')
// (19, 18, 'lutff_0/in_3')
// (19, 18, 'sp4_r_v_b_32')
// (19, 18, 'sp4_v_b_28')
// (19, 18, 'sp4_v_b_32')
// (19, 19, 'local_g1_5')
// (19, 19, 'lutff_3/in_3')
// (19, 19, 'sp4_r_v_b_21')
// (19, 19, 'sp4_v_b_17')
// (19, 19, 'sp4_v_b_21')
// (19, 20, 'sp4_r_v_b_8')
// (19, 20, 'sp4_v_b_4')
// (19, 20, 'sp4_v_b_8')
// (19, 21, 'sp4_r_v_b_45')
// (19, 22, 'sp4_r_v_b_32')
// (19, 23, 'sp4_r_v_b_21')
// (19, 24, 'sp4_r_v_b_8')
// (20, 8, 'sp4_v_t_44')
// (20, 9, 'sp4_v_b_44')
// (20, 10, 'sp4_v_b_33')
// (20, 11, 'local_g0_4')
// (20, 11, 'lutff_3/in_3')
// (20, 11, 'sp4_v_b_20')
// (20, 12, 'local_g0_3')
// (20, 12, 'lutff_4/in_3')
// (20, 12, 'sp12_h_r_11')
// (20, 12, 'sp4_h_l_38')
// (20, 12, 'sp4_h_r_29')
// (20, 12, 'sp4_h_r_7')
// (20, 12, 'sp4_v_b_9')
// (20, 12, 'sp4_v_t_45')
// (20, 13, 'sp4_v_b_45')
// (20, 14, 'sp4_v_b_32')
// (20, 15, 'sp4_v_b_21')
// (20, 16, 'local_g1_0')
// (20, 16, 'lutff_4/in_3')
// (20, 16, 'sp4_h_r_8')
// (20, 16, 'sp4_v_b_8')
// (20, 16, 'sp4_v_t_45')
// (20, 17, 'sp4_v_b_45')
// (20, 18, 'sp4_v_b_32')
// (20, 19, 'local_g0_5')
// (20, 19, 'lutff_4/in_3')
// (20, 19, 'sp4_v_b_21')
// (20, 20, 'local_g1_0')
// (20, 20, 'lutff_4/in_3')
// (20, 20, 'sp4_v_b_8')
// (20, 20, 'sp4_v_t_45')
// (20, 21, 'local_g3_5')
// (20, 21, 'lutff_3/in_3')
// (20, 21, 'sp4_v_b_45')
// (20, 22, 'sp4_v_b_32')
// (20, 23, 'sp4_v_b_21')
// (20, 24, 'sp4_v_b_8')
// (21, 9, 'sp4_r_v_b_40')
// (21, 10, 'sp4_r_v_b_29')
// (21, 11, 'local_g3_0')
// (21, 11, 'lutff_4/in_3')
// (21, 11, 'sp4_r_v_b_16')
// (21, 12, 'local_g0_4')
// (21, 12, 'lutff_4/in_0')
// (21, 12, 'sp12_h_r_12')
// (21, 12, 'sp4_h_r_18')
// (21, 12, 'sp4_h_r_40')
// (21, 12, 'sp4_r_v_b_5')
// (21, 13, 'sp4_r_v_b_47')
// (21, 14, 'sp4_r_v_b_34')
// (21, 15, 'local_g3_7')
// (21, 15, 'lutff_7/in_3')
// (21, 15, 'sp4_r_v_b_23')
// (21, 16, 'sp4_h_r_21')
// (21, 16, 'sp4_r_v_b_10')
// (21, 17, 'local_g2_4')
// (21, 17, 'lutff_3/in_3')
// (21, 17, 'sp4_r_v_b_36')
// (21, 18, 'sp4_r_v_b_25')
// (21, 19, 'sp4_r_v_b_12')
// (21, 20, 'local_g1_1')
// (21, 20, 'lutff_4/in_0')
// (21, 20, 'sp4_r_v_b_1')
// (21, 21, 'sp4_r_v_b_36')
// (21, 22, 'sp4_r_v_b_25')
// (21, 23, 'local_g2_4')
// (21, 23, 'lutff_2/in_0')
// (21, 23, 'sp4_r_v_b_12')
// (21, 24, 'local_g1_1')
// (21, 24, 'lutff_0/in_0')
// (21, 24, 'sp4_r_v_b_1')
// (22, 8, 'sp4_v_t_40')
// (22, 9, 'sp4_v_b_40')
// (22, 10, 'sp4_v_b_29')
// (22, 11, 'sp4_v_b_16')
// (22, 12, 'local_g1_7')
// (22, 12, 'lutff_4/in_0')
// (22, 12, 'sp12_h_r_15')
// (22, 12, 'sp4_h_l_40')
// (22, 12, 'sp4_h_r_31')
// (22, 12, 'sp4_v_b_5')
// (22, 12, 'sp4_v_t_47')
// (22, 13, 'local_g2_7')
// (22, 13, 'lutff_5/in_0')
// (22, 13, 'sp4_v_b_47')
// (22, 14, 'local_g3_2')
// (22, 14, 'lutff_4/in_3')
// (22, 14, 'sp4_v_b_34')
// (22, 15, 'sp4_v_b_23')
// (22, 16, 'sp4_h_r_32')
// (22, 16, 'sp4_v_b_10')
// (22, 16, 'sp4_v_t_36')
// (22, 17, 'sp4_v_b_36')
// (22, 18, 'sp4_v_b_25')
// (22, 19, 'local_g0_4')
// (22, 19, 'lutff_1/in_3')
// (22, 19, 'sp4_v_b_12')
// (22, 20, 'sp4_v_b_1')
// (22, 20, 'sp4_v_t_36')
// (22, 21, 'local_g3_4')
// (22, 21, 'lutff_4/in_3')
// (22, 21, 'sp4_v_b_36')
// (22, 22, 'sp4_v_b_25')
// (22, 23, 'local_g1_4')
// (22, 23, 'lutff_4/in_3')
// (22, 23, 'sp4_v_b_12')
// (22, 24, 'sp4_v_b_1')
// (23, 9, 'sp4_r_v_b_36')
// (23, 10, 'sp4_r_v_b_25')
// (23, 11, 'local_g2_4')
// (23, 11, 'lutff_1/in_3')
// (23, 11, 'sp4_r_v_b_12')
// (23, 12, 'local_g0_0')
// (23, 12, 'lutff_4/in_0')
// (23, 12, 'sp12_h_r_16')
// (23, 12, 'sp4_h_r_42')
// (23, 12, 'sp4_r_v_b_1')
// (23, 13, 'local_g3_2')
// (23, 13, 'lutff_1/in_0')
// (23, 13, 'sp4_r_v_b_42')
// (23, 14, 'local_g0_7')
// (23, 14, 'lutff_4/in_3')
// (23, 14, 'sp4_r_v_b_31')
// (23, 15, 'local_g3_2')
// (23, 15, 'lutff_4/in_3')
// (23, 15, 'sp4_r_v_b_18')
// (23, 16, 'local_g2_5')
// (23, 16, 'lutff_4/in_3')
// (23, 16, 'sp4_h_r_45')
// (23, 16, 'sp4_r_v_b_7')
// (23, 17, 'local_g2_6')
// (23, 17, 'lutff_5/in_3')
// (23, 17, 'sp4_r_v_b_38')
// (23, 18, 'local_g1_3')
// (23, 18, 'lutff_3/in_3')
// (23, 18, 'sp4_r_v_b_27')
// (23, 19, 'sp4_r_v_b_14')
// (23, 20, 'local_g1_3')
// (23, 20, 'lutff_4/in_0')
// (23, 20, 'sp4_r_v_b_3')
// (24, 8, 'sp4_v_t_36')
// (24, 9, 'sp4_v_b_36')
// (24, 10, 'sp4_v_b_25')
// (24, 11, 'sp4_v_b_12')
// (24, 12, 'sp12_h_r_19')
// (24, 12, 'sp4_h_l_42')
// (24, 12, 'sp4_v_b_1')
// (24, 12, 'sp4_v_t_42')
// (24, 13, 'sp4_v_b_42')
// (24, 14, 'local_g2_7')
// (24, 14, 'lutff_4/in_3')
// (24, 14, 'sp4_v_b_31')
// (24, 15, 'local_g1_2')
// (24, 15, 'lutff_2/in_3')
// (24, 15, 'sp4_v_b_18')
// (24, 16, 'sp4_h_l_45')
// (24, 16, 'sp4_v_b_7')
// (24, 16, 'sp4_v_t_38')
// (24, 17, 'local_g3_6')
// (24, 17, 'lutff_4/in_3')
// (24, 17, 'sp4_v_b_38')
// (24, 18, 'sp4_v_b_27')
// (24, 19, 'sp4_v_b_14')
// (24, 20, 'sp4_v_b_3')
// (25, 12, 'sp12_h_r_20')
// (26, 12, 'sp12_h_r_23')
// (27, 12, 'sp12_h_l_23')

reg n36 = 0;
// (3, 13, 'sp12_h_r_0')
// (4, 13, 'sp12_h_r_3')
// (5, 13, 'sp12_h_r_4')
// (6, 13, 'sp12_h_r_7')
// (7, 13, 'sp12_h_r_8')
// (8, 13, 'sp12_h_r_11')
// (9, 13, 'local_g0_4')
// (9, 13, 'lutff_1/in_3')
// (9, 13, 'sp12_h_r_12')
// (10, 13, 'sp12_h_r_15')
// (11, 13, 'sp12_h_r_16')
// (12, 12, 'local_g3_6')
// (12, 12, 'lutff_4/in_3')
// (12, 12, 'neigh_op_tnr_6')
// (12, 13, 'neigh_op_rgt_6')
// (12, 13, 'sp12_h_r_19')
// (12, 14, 'neigh_op_bnr_6')
// (13, 12, 'neigh_op_top_6')
// (13, 13, 'lutff_6/out')
// (13, 13, 'sp12_h_r_20')
// (13, 14, 'neigh_op_bot_6')
// (14, 12, 'neigh_op_tnl_6')
// (14, 13, 'neigh_op_lft_6')
// (14, 13, 'sp12_h_r_23')
// (14, 14, 'neigh_op_bnl_6')
// (15, 13, 'sp12_h_l_23')

reg n37 = 0;
// (3, 18, 'sp12_h_r_0')
// (4, 18, 'sp12_h_r_3')
// (5, 18, 'sp12_h_r_4')
// (6, 18, 'sp12_h_r_7')
// (7, 18, 'sp12_h_r_8')
// (8, 17, 'neigh_op_tnr_2')
// (8, 18, 'neigh_op_rgt_2')
// (8, 18, 'sp12_h_r_11')
// (8, 19, 'neigh_op_bnr_2')
// (9, 17, 'neigh_op_top_2')
// (9, 18, 'lutff_2/out')
// (9, 18, 'sp12_h_r_12')
// (9, 19, 'neigh_op_bot_2')
// (10, 17, 'neigh_op_tnl_2')
// (10, 18, 'neigh_op_lft_2')
// (10, 18, 'sp12_h_r_15')
// (10, 19, 'neigh_op_bnl_2')
// (11, 18, 'sp12_h_r_16')
// (12, 18, 'sp12_h_r_19')
// (13, 18, 'local_g1_4')
// (13, 18, 'lutff_6/in_1')
// (13, 18, 'sp12_h_r_20')
// (14, 18, 'sp12_h_r_23')
// (15, 18, 'sp12_h_l_23')

wire io_4_33_0;
// (3, 32, 'neigh_op_tnr_0')
// (3, 32, 'neigh_op_tnr_4')
// (4, 29, 'sp12_h_r_0')
// (4, 29, 'sp12_v_t_23')
// (4, 30, 'sp12_v_b_23')
// (4, 31, 'sp12_v_b_20')
// (4, 32, 'neigh_op_top_0')
// (4, 32, 'neigh_op_top_4')
// (4, 32, 'sp12_v_b_19')
// (4, 33, 'io_0/D_IN_0')
// (4, 33, 'io_0/PAD')
// (4, 33, 'span12_vert_16')
// (5, 29, 'sp12_h_r_3')
// (5, 32, 'neigh_op_tnl_0')
// (5, 32, 'neigh_op_tnl_4')
// (6, 29, 'sp12_h_r_4')
// (7, 29, 'sp12_h_r_7')
// (8, 29, 'sp12_h_r_8')
// (9, 29, 'sp12_h_r_11')
// (10, 29, 'sp12_h_r_12')
// (11, 29, 'sp12_h_r_15')
// (12, 29, 'sp12_h_r_16')
// (13, 29, 'sp12_h_r_19')
// (14, 29, 'sp12_h_r_20')
// (15, 29, 'sp12_h_r_23')
// (16, 17, 'sp12_v_t_23')
// (16, 18, 'sp12_v_b_23')
// (16, 19, 'sp12_v_b_20')
// (16, 20, 'sp12_v_b_19')
// (16, 21, 'sp12_v_b_16')
// (16, 22, 'sp12_v_b_15')
// (16, 23, 'sp12_v_b_12')
// (16, 24, 'local_g3_3')
// (16, 24, 'lutff_5/in_3')
// (16, 24, 'sp12_v_b_11')
// (16, 25, 'sp12_v_b_8')
// (16, 26, 'sp12_v_b_7')
// (16, 27, 'sp12_v_b_4')
// (16, 28, 'sp12_v_b_3')
// (16, 29, 'sp12_h_l_23')
// (16, 29, 'sp12_v_b_0')

wire io_4_33_1;
// (3, 32, 'neigh_op_tnr_2')
// (3, 32, 'neigh_op_tnr_6')
// (4, 23, 'sp12_h_r_0')
// (4, 23, 'sp12_v_t_23')
// (4, 24, 'sp12_v_b_23')
// (4, 25, 'sp12_v_b_20')
// (4, 26, 'sp12_v_b_19')
// (4, 27, 'sp12_v_b_16')
// (4, 28, 'sp12_v_b_15')
// (4, 29, 'sp12_v_b_12')
// (4, 30, 'sp12_v_b_11')
// (4, 31, 'sp12_v_b_8')
// (4, 32, 'neigh_op_top_2')
// (4, 32, 'neigh_op_top_6')
// (4, 32, 'sp12_v_b_7')
// (4, 33, 'io_1/D_IN_0')
// (4, 33, 'io_1/PAD')
// (4, 33, 'span12_vert_4')
// (5, 23, 'sp12_h_r_3')
// (5, 32, 'neigh_op_tnl_2')
// (5, 32, 'neigh_op_tnl_6')
// (6, 23, 'sp12_h_r_4')
// (7, 23, 'sp12_h_r_7')
// (8, 23, 'sp12_h_r_8')
// (9, 23, 'sp12_h_r_11')
// (10, 23, 'sp12_h_r_12')
// (11, 23, 'sp12_h_r_15')
// (12, 23, 'sp12_h_r_16')
// (13, 23, 'sp12_h_r_19')
// (14, 23, 'sp12_h_r_20')
// (15, 23, 'sp12_h_r_23')
// (16, 23, 'sp12_h_l_23')
// (16, 23, 'sp12_v_t_23')
// (16, 24, 'local_g2_7')
// (16, 24, 'lutff_4/in_3')
// (16, 24, 'sp12_v_b_23')
// (16, 25, 'sp12_v_b_20')
// (16, 26, 'sp12_v_b_19')
// (16, 27, 'sp12_v_b_16')
// (16, 28, 'sp12_v_b_15')
// (16, 29, 'sp12_v_b_12')
// (16, 30, 'sp12_v_b_11')
// (16, 31, 'sp12_v_b_8')
// (16, 32, 'sp12_v_b_7')
// (16, 33, 'span12_vert_4')

reg io_4_0_0 = 0;
// (4, 0, 'io_0/D_OUT_0')
// (4, 0, 'io_0/PAD')
// (4, 0, 'local_g0_2')
// (4, 0, 'span12_vert_18')
// (4, 1, 'sp12_v_b_18')
// (4, 2, 'sp12_v_b_17')
// (4, 3, 'sp12_v_b_14')
// (4, 4, 'sp12_v_b_13')
// (4, 5, 'sp12_v_b_10')
// (4, 6, 'sp12_v_b_9')
// (4, 7, 'sp12_v_b_6')
// (4, 8, 'sp12_v_b_5')
// (4, 9, 'sp12_v_b_2')
// (4, 10, 'sp12_h_r_1')
// (4, 10, 'sp12_v_b_1')
// (5, 10, 'sp12_h_r_2')
// (6, 9, 'neigh_op_tnr_7')
// (6, 10, 'neigh_op_rgt_7')
// (6, 10, 'sp12_h_r_5')
// (6, 10, 'sp4_h_r_3')
// (6, 11, 'neigh_op_bnr_7')
// (7, 9, 'neigh_op_top_7')
// (7, 10, 'lutff_7/out')
// (7, 10, 'sp12_h_r_6')
// (7, 10, 'sp4_h_r_14')
// (7, 11, 'neigh_op_bot_7')
// (8, 9, 'neigh_op_tnl_7')
// (8, 10, 'neigh_op_lft_7')
// (8, 10, 'sp12_h_r_9')
// (8, 10, 'sp4_h_r_27')
// (8, 11, 'neigh_op_bnl_7')
// (9, 10, 'local_g2_6')
// (9, 10, 'lutff_3/in_3')
// (9, 10, 'sp12_h_r_10')
// (9, 10, 'sp4_h_r_38')
// (10, 10, 'sp12_h_r_13')
// (10, 10, 'sp4_h_l_38')
// (11, 10, 'sp12_h_r_14')
// (12, 10, 'sp12_h_r_17')
// (13, 10, 'sp12_h_r_18')
// (14, 10, 'sp12_h_r_21')
// (15, 10, 'sp12_h_r_22')
// (16, 10, 'sp12_h_l_22')

reg n41 = 0;
// (4, 10, 'sp12_h_r_0')
// (5, 10, 'sp12_h_r_3')
// (6, 10, 'sp12_h_r_4')
// (7, 10, 'local_g0_7')
// (7, 10, 'lutff_6/in_3')
// (7, 10, 'sp12_h_r_7')
// (8, 10, 'sp12_h_r_8')
// (9, 10, 'sp12_h_r_11')
// (10, 10, 'sp12_h_r_12')
// (11, 10, 'sp12_h_r_15')
// (12, 10, 'sp12_h_r_16')
// (13, 10, 'sp12_h_r_19')
// (14, 10, 'sp12_h_r_20')
// (15, 10, 'local_g1_5')
// (15, 10, 'lutff_5/in_3')
// (15, 10, 'sp12_h_r_23')
// (15, 10, 'sp4_h_r_5')
// (16, 10, 'sp12_h_l_23')
// (16, 10, 'sp12_h_r_0')
// (16, 10, 'sp4_h_r_16')
// (17, 10, 'sp12_h_r_3')
// (17, 10, 'sp4_h_r_29')
// (18, 10, 'sp12_h_r_4')
// (18, 10, 'sp4_h_r_40')
// (19, 9, 'neigh_op_tnr_0')
// (19, 10, 'neigh_op_rgt_0')
// (19, 10, 'sp12_h_r_7')
// (19, 10, 'sp4_h_l_40')
// (19, 10, 'sp4_h_r_5')
// (19, 11, 'neigh_op_bnr_0')
// (20, 9, 'neigh_op_top_0')
// (20, 10, 'local_g0_0')
// (20, 10, 'lutff_0/in_2')
// (20, 10, 'lutff_0/out')
// (20, 10, 'sp12_h_r_8')
// (20, 10, 'sp4_h_r_16')
// (20, 11, 'neigh_op_bot_0')
// (21, 9, 'neigh_op_tnl_0')
// (21, 10, 'neigh_op_lft_0')
// (21, 10, 'sp12_h_r_11')
// (21, 10, 'sp4_h_r_29')
// (21, 11, 'neigh_op_bnl_0')
// (22, 10, 'sp12_h_r_12')
// (22, 10, 'sp4_h_r_40')
// (23, 10, 'sp12_h_r_15')
// (23, 10, 'sp4_h_l_40')
// (24, 10, 'sp12_h_r_16')
// (25, 10, 'sp12_h_r_19')
// (26, 10, 'sp12_h_r_20')
// (27, 10, 'sp12_h_r_23')
// (28, 10, 'sp12_h_l_23')

reg n42 = 0;
// (4, 12, 'sp12_h_r_1')
// (5, 12, 'sp12_h_r_2')
// (6, 12, 'sp12_h_r_5')
// (7, 12, 'sp12_h_r_6')
// (8, 12, 'sp12_h_r_9')
// (9, 12, 'sp12_h_r_10')
// (9, 13, 'sp4_r_v_b_40')
// (9, 14, 'sp4_r_v_b_29')
// (9, 15, 'sp4_r_v_b_16')
// (9, 16, 'local_g1_5')
// (9, 16, 'lutff_7/in_1')
// (9, 16, 'sp4_r_v_b_5')
// (9, 17, 'local_g2_4')
// (9, 17, 'lutff_7/in_3')
// (9, 17, 'sp4_r_v_b_36')
// (9, 18, 'sp4_r_v_b_25')
// (9, 19, 'sp4_r_v_b_12')
// (9, 20, 'sp4_r_v_b_1')
// (10, 11, 'neigh_op_tnr_3')
// (10, 12, 'neigh_op_rgt_3')
// (10, 12, 'sp12_h_r_13')
// (10, 12, 'sp4_h_r_11')
// (10, 12, 'sp4_v_t_40')
// (10, 13, 'neigh_op_bnr_3')
// (10, 13, 'sp4_v_b_40')
// (10, 14, 'sp4_v_b_29')
// (10, 15, 'sp4_v_b_16')
// (10, 16, 'sp4_v_b_5')
// (10, 16, 'sp4_v_t_36')
// (10, 17, 'sp4_v_b_36')
// (10, 18, 'sp4_v_b_25')
// (10, 19, 'local_g0_4')
// (10, 19, 'lutff_3/in_3')
// (10, 19, 'sp4_r_v_b_38')
// (10, 19, 'sp4_v_b_12')
// (10, 20, 'local_g1_1')
// (10, 20, 'lutff_1/in_3')
// (10, 20, 'sp4_r_v_b_27')
// (10, 20, 'sp4_v_b_1')
// (10, 21, 'sp4_r_v_b_14')
// (10, 22, 'sp4_r_v_b_3')
// (11, 3, 'sp12_v_t_22')
// (11, 4, 'sp12_v_b_22')
// (11, 5, 'sp12_v_b_21')
// (11, 6, 'sp12_v_b_18')
// (11, 7, 'sp12_v_b_17')
// (11, 8, 'sp12_v_b_14')
// (11, 9, 'sp12_v_b_13')
// (11, 10, 'sp12_v_b_10')
// (11, 11, 'neigh_op_top_3')
// (11, 11, 'sp12_h_r_1')
// (11, 11, 'sp12_v_b_9')
// (11, 11, 'sp12_v_t_22')
// (11, 12, 'lutff_3/out')
// (11, 12, 'sp12_h_r_14')
// (11, 12, 'sp12_v_b_22')
// (11, 12, 'sp12_v_b_6')
// (11, 12, 'sp4_h_r_22')
// (11, 12, 'sp4_r_v_b_39')
// (11, 13, 'local_g1_3')
// (11, 13, 'lutff_1/in_3')
// (11, 13, 'neigh_op_bot_3')
// (11, 13, 'sp12_v_b_21')
// (11, 13, 'sp12_v_b_5')
// (11, 13, 'sp4_r_v_b_26')
// (11, 14, 'sp12_v_b_18')
// (11, 14, 'sp12_v_b_2')
// (11, 14, 'sp4_r_v_b_15')
// (11, 15, 'sp12_h_r_1')
// (11, 15, 'sp12_v_b_1')
// (11, 15, 'sp12_v_b_17')
// (11, 15, 'sp4_r_v_b_2')
// (11, 16, 'sp12_v_b_14')
// (11, 16, 'sp4_r_v_b_40')
// (11, 17, 'sp12_v_b_13')
// (11, 17, 'sp4_r_v_b_29')
// (11, 18, 'sp12_v_b_10')
// (11, 18, 'sp4_r_v_b_16')
// (11, 18, 'sp4_v_t_38')
// (11, 19, 'sp12_v_b_9')
// (11, 19, 'sp4_r_v_b_5')
// (11, 19, 'sp4_v_b_38')
// (11, 20, 'sp12_v_b_6')
// (11, 20, 'sp4_r_v_b_36')
// (11, 20, 'sp4_v_b_27')
// (11, 21, 'sp12_v_b_5')
// (11, 21, 'sp4_r_v_b_25')
// (11, 21, 'sp4_v_b_14')
// (11, 22, 'local_g2_2')
// (11, 22, 'lutff_7/in_3')
// (11, 22, 'sp12_v_b_2')
// (11, 22, 'sp4_h_r_3')
// (11, 22, 'sp4_r_v_b_12')
// (11, 22, 'sp4_v_b_3')
// (11, 23, 'sp12_h_r_1')
// (11, 23, 'sp12_v_b_1')
// (11, 23, 'sp4_r_v_b_1')
// (12, 11, 'neigh_op_tnl_3')
// (12, 11, 'sp12_h_r_2')
// (12, 11, 'sp4_v_t_39')
// (12, 12, 'neigh_op_lft_3')
// (12, 12, 'sp12_h_r_17')
// (12, 12, 'sp4_h_r_35')
// (12, 12, 'sp4_v_b_39')
// (12, 13, 'local_g3_3')
// (12, 13, 'lutff_3/in_3')
// (12, 13, 'neigh_op_bnl_3')
// (12, 13, 'sp4_v_b_26')
// (12, 14, 'sp4_v_b_15')
// (12, 15, 'sp12_h_r_2')
// (12, 15, 'sp4_h_r_8')
// (12, 15, 'sp4_v_b_2')
// (12, 15, 'sp4_v_t_40')
// (12, 16, 'sp4_v_b_40')
// (12, 17, 'sp4_v_b_29')
// (12, 18, 'sp4_v_b_16')
// (12, 19, 'local_g1_5')
// (12, 19, 'lutff_3/in_3')
// (12, 19, 'sp4_v_b_5')
// (12, 19, 'sp4_v_t_36')
// (12, 20, 'local_g2_4')
// (12, 20, 'lutff_3/in_3')
// (12, 20, 'sp4_v_b_36')
// (12, 21, 'sp4_v_b_25')
// (12, 22, 'sp4_h_r_14')
// (12, 22, 'sp4_v_b_12')
// (12, 23, 'sp12_h_r_2')
// (12, 23, 'sp4_v_b_1')
// (13, 11, 'sp12_h_r_5')
// (13, 12, 'sp12_h_r_18')
// (13, 12, 'sp4_h_r_46')
// (13, 13, 'sp4_r_v_b_46')
// (13, 14, 'local_g2_3')
// (13, 14, 'lutff_4/in_3')
// (13, 14, 'sp4_r_v_b_35')
// (13, 15, 'sp12_h_r_5')
// (13, 15, 'sp4_h_r_21')
// (13, 15, 'sp4_r_v_b_22')
// (13, 16, 'local_g2_3')
// (13, 16, 'lutff_1/in_0')
// (13, 16, 'sp4_r_v_b_11')
// (13, 22, 'sp4_h_r_27')
// (13, 23, 'sp12_h_r_5')
// (14, 11, 'sp12_h_r_6')
// (14, 12, 'sp12_h_r_21')
// (14, 12, 'sp4_h_l_46')
// (14, 12, 'sp4_v_t_46')
// (14, 13, 'local_g2_6')
// (14, 13, 'lutff_3/in_3')
// (14, 13, 'sp4_v_b_46')
// (14, 14, 'sp4_v_b_35')
// (14, 15, 'sp12_h_r_6')
// (14, 15, 'sp4_h_r_32')
// (14, 15, 'sp4_v_b_22')
// (14, 16, 'sp4_h_r_5')
// (14, 16, 'sp4_v_b_11')
// (14, 22, 'local_g3_6')
// (14, 22, 'lutff_2/in_3')
// (14, 22, 'sp4_h_r_38')
// (14, 23, 'sp12_h_r_6')
// (15, 11, 'sp12_h_r_9')
// (15, 12, 'sp12_h_r_22')
// (15, 15, 'local_g3_5')
// (15, 15, 'lutff_3/in_3')
// (15, 15, 'sp12_h_r_9')
// (15, 15, 'sp4_h_r_45')
// (15, 16, 'sp4_h_r_16')
// (15, 16, 'sp4_r_v_b_45')
// (15, 17, 'local_g2_0')
// (15, 17, 'lutff_3/in_3')
// (15, 17, 'sp4_r_v_b_32')
// (15, 18, 'local_g3_5')
// (15, 18, 'lutff_3/in_3')
// (15, 18, 'sp4_r_v_b_21')
// (15, 19, 'local_g2_0')
// (15, 19, 'lutff_3/in_3')
// (15, 19, 'sp4_r_v_b_8')
// (15, 22, 'sp4_h_l_38')
// (15, 23, 'sp12_h_r_9')
// (16, 0, 'span12_vert_22')
// (16, 1, 'sp12_v_b_22')
// (16, 2, 'sp12_v_b_21')
// (16, 3, 'sp12_v_b_18')
// (16, 4, 'sp12_v_b_17')
// (16, 5, 'sp12_v_b_14')
// (16, 6, 'sp12_v_b_13')
// (16, 7, 'sp12_v_b_10')
// (16, 8, 'sp12_v_b_9')
// (16, 9, 'sp12_v_b_6')
// (16, 10, 'sp12_v_b_5')
// (16, 11, 'local_g3_2')
// (16, 11, 'lutff_3/in_0')
// (16, 11, 'sp12_h_r_10')
// (16, 11, 'sp12_v_b_2')
// (16, 12, 'sp12_h_l_22')
// (16, 12, 'sp12_h_r_1')
// (16, 12, 'sp12_v_b_1')
// (16, 12, 'sp12_v_t_22')
// (16, 13, 'local_g2_6')
// (16, 13, 'lutff_3/in_1')
// (16, 13, 'sp12_v_b_22')
// (16, 14, 'sp12_v_b_21')
// (16, 15, 'sp12_h_r_10')
// (16, 15, 'sp12_v_b_18')
// (16, 15, 'sp4_h_l_45')
// (16, 15, 'sp4_v_t_45')
// (16, 16, 'local_g3_1')
// (16, 16, 'lutff_3/in_3')
// (16, 16, 'sp12_v_b_17')
// (16, 16, 'sp4_h_r_29')
// (16, 16, 'sp4_v_b_45')
// (16, 17, 'local_g3_6')
// (16, 17, 'lutff_3/in_0')
// (16, 17, 'sp12_v_b_14')
// (16, 17, 'sp4_v_b_32')
// (16, 18, 'local_g3_5')
// (16, 18, 'lutff_3/in_3')
// (16, 18, 'sp12_v_b_13')
// (16, 18, 'sp4_v_b_21')
// (16, 19, 'local_g0_0')
// (16, 19, 'lutff_1/in_1')
// (16, 19, 'sp12_v_b_10')
// (16, 19, 'sp4_h_r_2')
// (16, 19, 'sp4_v_b_8')
// (16, 20, 'sp12_v_b_9')
// (16, 21, 'local_g2_6')
// (16, 21, 'lutff_1/in_3')
// (16, 21, 'sp12_v_b_6')
// (16, 22, 'sp12_v_b_5')
// (16, 23, 'sp12_h_r_10')
// (16, 23, 'sp12_v_b_2')
// (16, 24, 'sp12_h_r_1')
// (16, 24, 'sp12_v_b_1')
// (17, 11, 'sp12_h_r_13')
// (17, 12, 'sp12_h_r_2')
// (17, 15, 'sp12_h_r_13')
// (17, 15, 'sp4_h_r_6')
// (17, 16, 'sp4_h_r_40')
// (17, 19, 'sp4_h_r_15')
// (17, 23, 'sp12_h_r_13')
// (17, 24, 'sp12_h_r_2')
// (18, 11, 'sp12_h_r_14')
// (18, 12, 'local_g1_5')
// (18, 12, 'lutff_3/in_3')
// (18, 12, 'sp12_h_r_5')
// (18, 15, 'sp12_h_r_14')
// (18, 15, 'sp4_h_r_19')
// (18, 16, 'sp4_h_l_40')
// (18, 16, 'sp4_h_r_1')
// (18, 19, 'sp4_h_r_26')
// (18, 23, 'sp12_h_r_14')
// (18, 24, 'sp12_h_r_5')
// (19, 11, 'local_g1_1')
// (19, 11, 'lutff_3/in_3')
// (19, 11, 'sp12_h_r_17')
// (19, 11, 'sp4_h_r_8')
// (19, 12, 'sp12_h_r_6')
// (19, 15, 'sp12_h_r_17')
// (19, 15, 'sp4_h_r_30')
// (19, 16, 'local_g0_4')
// (19, 16, 'lutff_3/in_3')
// (19, 16, 'sp4_h_r_12')
// (19, 19, 'local_g2_7')
// (19, 19, 'lutff_2/in_3')
// (19, 19, 'sp4_h_r_39')
// (19, 20, 'sp4_r_v_b_39')
// (19, 21, 'sp4_r_v_b_26')
// (19, 22, 'sp4_r_v_b_15')
// (19, 23, 'sp12_h_r_17')
// (19, 23, 'sp4_r_v_b_2')
// (19, 24, 'sp12_h_r_6')
// (19, 24, 'sp4_r_v_b_40')
// (19, 25, 'sp4_r_v_b_29')
// (19, 26, 'sp4_r_v_b_16')
// (19, 27, 'sp4_r_v_b_5')
// (20, 11, 'local_g1_2')
// (20, 11, 'lutff_2/in_3')
// (20, 11, 'sp12_h_r_18')
// (20, 11, 'sp4_h_r_21')
// (20, 12, 'local_g1_1')
// (20, 12, 'lutff_3/in_3')
// (20, 12, 'sp12_h_r_9')
// (20, 15, 'sp12_h_r_18')
// (20, 15, 'sp4_h_r_43')
// (20, 16, 'local_g3_1')
// (20, 16, 'lutff_3/in_3')
// (20, 16, 'sp4_h_r_25')
// (20, 16, 'sp4_r_v_b_43')
// (20, 17, 'local_g0_6')
// (20, 17, 'lutff_7/in_3')
// (20, 17, 'sp4_r_v_b_30')
// (20, 18, 'sp4_r_v_b_19')
// (20, 19, 'local_g1_6')
// (20, 19, 'lutff_3/in_0')
// (20, 19, 'sp4_h_l_39')
// (20, 19, 'sp4_r_v_b_6')
// (20, 19, 'sp4_v_t_39')
// (20, 20, 'local_g3_7')
// (20, 20, 'lutff_3/in_3')
// (20, 20, 'sp4_v_b_39')
// (20, 21, 'local_g2_2')
// (20, 21, 'lutff_1/in_3')
// (20, 21, 'sp4_v_b_26')
// (20, 22, 'sp4_v_b_15')
// (20, 23, 'local_g0_2')
// (20, 23, 'lutff_6/in_0')
// (20, 23, 'sp12_h_r_18')
// (20, 23, 'sp4_v_b_2')
// (20, 23, 'sp4_v_t_40')
// (20, 24, 'sp12_h_r_9')
// (20, 24, 'sp4_v_b_40')
// (20, 25, 'local_g3_5')
// (20, 25, 'lutff_3/in_3')
// (20, 25, 'sp4_v_b_29')
// (20, 26, 'sp4_v_b_16')
// (20, 27, 'sp4_v_b_5')
// (21, 11, 'local_g1_5')
// (21, 11, 'lutff_3/in_3')
// (21, 11, 'sp12_h_r_21')
// (21, 11, 'sp4_h_r_32')
// (21, 12, 'local_g0_2')
// (21, 12, 'lutff_3/in_3')
// (21, 12, 'sp12_h_r_10')
// (21, 13, 'sp4_r_v_b_42')
// (21, 14, 'sp4_r_v_b_31')
// (21, 15, 'local_g0_5')
// (21, 15, 'lutff_5/in_0')
// (21, 15, 'sp12_h_r_21')
// (21, 15, 'sp4_h_l_43')
// (21, 15, 'sp4_h_r_10')
// (21, 15, 'sp4_r_v_b_18')
// (21, 15, 'sp4_v_t_43')
// (21, 16, 'sp4_h_r_36')
// (21, 16, 'sp4_r_v_b_7')
// (21, 16, 'sp4_v_b_43')
// (21, 17, 'local_g2_6')
// (21, 17, 'lutff_1/in_3')
// (21, 17, 'sp4_r_v_b_42')
// (21, 17, 'sp4_v_b_30')
// (21, 18, 'local_g1_3')
// (21, 18, 'lutff_5/in_3')
// (21, 18, 'sp4_r_v_b_31')
// (21, 18, 'sp4_v_b_19')
// (21, 19, 'sp4_r_v_b_18')
// (21, 19, 'sp4_v_b_6')
// (21, 20, 'local_g1_7')
// (21, 20, 'lutff_3/in_3')
// (21, 20, 'sp4_r_v_b_7')
// (21, 23, 'sp12_h_r_21')
// (21, 24, 'sp12_h_r_10')
// (22, 11, 'sp12_h_r_22')
// (22, 11, 'sp4_h_r_45')
// (22, 12, 'local_g1_5')
// (22, 12, 'lutff_3/in_3')
// (22, 12, 'sp12_h_r_13')
// (22, 12, 'sp4_r_v_b_36')
// (22, 12, 'sp4_v_t_42')
// (22, 13, 'local_g0_1')
// (22, 13, 'lutff_2/in_1')
// (22, 13, 'sp4_r_v_b_25')
// (22, 13, 'sp4_v_b_42')
// (22, 14, 'local_g2_4')
// (22, 14, 'lutff_3/in_3')
// (22, 14, 'sp4_r_v_b_12')
// (22, 14, 'sp4_v_b_31')
// (22, 15, 'sp12_h_r_22')
// (22, 15, 'sp4_h_r_23')
// (22, 15, 'sp4_r_v_b_1')
// (22, 15, 'sp4_v_b_18')
// (22, 16, 'local_g0_7')
// (22, 16, 'lutff_0/in_3')
// (22, 16, 'sp4_h_l_36')
// (22, 16, 'sp4_v_b_7')
// (22, 16, 'sp4_v_t_42')
// (22, 17, 'sp4_v_b_42')
// (22, 18, 'sp4_v_b_31')
// (22, 19, 'sp4_r_v_b_38')
// (22, 19, 'sp4_v_b_18')
// (22, 20, 'sp4_r_v_b_27')
// (22, 20, 'sp4_v_b_7')
// (22, 21, 'local_g2_6')
// (22, 21, 'lutff_3/in_3')
// (22, 21, 'sp4_r_v_b_14')
// (22, 22, 'sp4_r_v_b_3')
// (22, 23, 'local_g0_6')
// (22, 23, 'lutff_3/in_3')
// (22, 23, 'sp12_h_r_22')
// (22, 24, 'local_g0_5')
// (22, 24, 'lutff_0/in_3')
// (22, 24, 'sp12_h_r_13')
// (23, 11, 'sp12_h_l_22')
// (23, 11, 'sp12_v_t_22')
// (23, 11, 'sp4_h_l_45')
// (23, 11, 'sp4_v_t_36')
// (23, 12, 'local_g0_6')
// (23, 12, 'lutff_3/in_3')
// (23, 12, 'sp12_h_r_14')
// (23, 12, 'sp12_v_b_22')
// (23, 12, 'sp4_v_b_36')
// (23, 13, 'sp12_v_b_21')
// (23, 13, 'sp4_v_b_25')
// (23, 14, 'local_g0_4')
// (23, 14, 'lutff_3/in_3')
// (23, 14, 'sp12_v_b_18')
// (23, 14, 'sp4_v_b_12')
// (23, 15, 'local_g1_1')
// (23, 15, 'lutff_3/in_3')
// (23, 15, 'sp12_h_l_22')
// (23, 15, 'sp12_v_b_17')
// (23, 15, 'sp4_h_r_34')
// (23, 15, 'sp4_v_b_1')
// (23, 16, 'local_g3_6')
// (23, 16, 'lutff_3/in_0')
// (23, 16, 'sp12_v_b_14')
// (23, 17, 'local_g3_5')
// (23, 17, 'lutff_0/in_0')
// (23, 17, 'sp12_v_b_13')
// (23, 18, 'local_g3_2')
// (23, 18, 'lutff_2/in_3')
// (23, 18, 'sp12_v_b_10')
// (23, 18, 'sp4_v_t_38')
// (23, 19, 'sp12_v_b_9')
// (23, 19, 'sp4_v_b_38')
// (23, 20, 'local_g2_6')
// (23, 20, 'lutff_3/in_3')
// (23, 20, 'sp12_v_b_6')
// (23, 20, 'sp4_v_b_27')
// (23, 21, 'sp12_v_b_5')
// (23, 21, 'sp4_v_b_14')
// (23, 22, 'sp12_v_b_2')
// (23, 22, 'sp4_v_b_3')
// (23, 23, 'sp12_h_l_22')
// (23, 23, 'sp12_v_b_1')
// (23, 24, 'sp12_h_r_14')
// (24, 12, 'sp12_h_r_17')
// (24, 12, 'sp4_r_v_b_41')
// (24, 13, 'sp4_r_v_b_28')
// (24, 14, 'local_g3_1')
// (24, 14, 'lutff_3/in_3')
// (24, 14, 'sp4_r_v_b_17')
// (24, 15, 'sp4_h_r_47')
// (24, 15, 'sp4_r_v_b_4')
// (24, 16, 'sp4_r_v_b_47')
// (24, 17, 'local_g0_1')
// (24, 17, 'lutff_3/in_0')
// (24, 17, 'sp4_r_v_b_34')
// (24, 18, 'sp4_r_v_b_23')
// (24, 19, 'sp4_r_v_b_10')
// (24, 24, 'sp12_h_r_17')
// (25, 11, 'sp4_v_t_41')
// (25, 12, 'sp12_h_r_18')
// (25, 12, 'sp4_v_b_41')
// (25, 13, 'sp4_v_b_28')
// (25, 14, 'sp4_v_b_17')
// (25, 15, 'sp4_h_l_47')
// (25, 15, 'sp4_v_b_4')
// (25, 15, 'sp4_v_t_47')
// (25, 16, 'sp4_v_b_47')
// (25, 17, 'sp4_v_b_34')
// (25, 18, 'sp4_v_b_23')
// (25, 19, 'sp4_v_b_10')
// (25, 24, 'sp12_h_r_18')
// (26, 12, 'sp12_h_r_21')
// (26, 24, 'sp12_h_r_21')
// (27, 12, 'sp12_h_r_22')
// (27, 24, 'sp12_h_r_22')
// (28, 12, 'sp12_h_l_22')
// (28, 24, 'sp12_h_l_22')

reg n43 = 0;
// (4, 12, 'sp4_h_r_2')
// (5, 12, 'sp4_h_r_15')
// (6, 12, 'sp4_h_r_26')
// (7, 12, 'local_g3_7')
// (7, 12, 'lutff_5/in_3')
// (7, 12, 'sp4_h_r_39')
// (8, 11, 'neigh_op_tnr_3')
// (8, 12, 'neigh_op_rgt_3')
// (8, 12, 'sp4_h_l_39')
// (8, 12, 'sp4_h_r_11')
// (8, 13, 'neigh_op_bnr_3')
// (9, 11, 'neigh_op_top_3')
// (9, 12, 'local_g0_6')
// (9, 12, 'lutff_3/in_1')
// (9, 12, 'lutff_3/out')
// (9, 12, 'sp4_h_r_22')
// (9, 13, 'neigh_op_bot_3')
// (10, 11, 'neigh_op_tnl_3')
// (10, 12, 'local_g1_3')
// (10, 12, 'lutff_1/in_3')
// (10, 12, 'neigh_op_lft_3')
// (10, 12, 'sp4_h_r_35')
// (10, 13, 'neigh_op_bnl_3')
// (11, 12, 'sp4_h_r_46')
// (12, 12, 'sp4_h_l_46')

reg n44 = 0;
// (4, 13, 'sp12_h_r_1')
// (5, 13, 'sp12_h_r_2')
// (6, 13, 'sp12_h_r_5')
// (7, 13, 'sp12_h_r_6')
// (8, 12, 'neigh_op_tnr_1')
// (8, 12, 'sp4_r_v_b_47')
// (8, 13, 'neigh_op_rgt_1')
// (8, 13, 'sp12_h_r_9')
// (8, 13, 'sp4_r_v_b_34')
// (8, 14, 'neigh_op_bnr_1')
// (8, 14, 'sp4_r_v_b_23')
// (8, 15, 'sp4_r_v_b_10')
// (8, 20, 'sp4_h_r_1')
// (9, 11, 'sp4_v_t_47')
// (9, 12, 'neigh_op_top_1')
// (9, 12, 'sp4_r_v_b_46')
// (9, 12, 'sp4_v_b_47')
// (9, 13, 'lutff_1/out')
// (9, 13, 'sp12_h_r_10')
// (9, 13, 'sp4_r_v_b_35')
// (9, 13, 'sp4_v_b_34')
// (9, 14, 'neigh_op_bot_1')
// (9, 14, 'sp4_r_v_b_22')
// (9, 14, 'sp4_v_b_23')
// (9, 15, 'local_g1_2')
// (9, 15, 'lutff_6/in_1')
// (9, 15, 'sp4_h_r_4')
// (9, 15, 'sp4_r_v_b_11')
// (9, 15, 'sp4_v_b_10')
// (9, 16, 'sp4_r_v_b_46')
// (9, 17, 'local_g2_3')
// (9, 17, 'lutff_6/in_3')
// (9, 17, 'sp4_r_v_b_35')
// (9, 18, 'sp4_r_v_b_22')
// (9, 19, 'sp4_r_v_b_11')
// (9, 20, 'sp4_h_r_12')
// (10, 11, 'sp4_v_t_46')
// (10, 12, 'neigh_op_tnl_1')
// (10, 12, 'sp4_v_b_46')
// (10, 13, 'neigh_op_lft_1')
// (10, 13, 'sp12_h_r_13')
// (10, 13, 'sp4_h_r_6')
// (10, 13, 'sp4_v_b_35')
// (10, 14, 'neigh_op_bnl_1')
// (10, 14, 'sp4_v_b_22')
// (10, 15, 'sp4_h_r_17')
// (10, 15, 'sp4_v_b_11')
// (10, 15, 'sp4_v_t_46')
// (10, 16, 'sp4_v_b_46')
// (10, 17, 'sp4_v_b_35')
// (10, 18, 'sp4_v_b_22')
// (10, 19, 'local_g0_3')
// (10, 19, 'lutff_2/in_3')
// (10, 19, 'sp4_v_b_11')
// (10, 20, 'local_g2_1')
// (10, 20, 'lutff_0/in_3')
// (10, 20, 'sp4_h_r_25')
// (11, 13, 'local_g0_3')
// (11, 13, 'lutff_0/in_3')
// (11, 13, 'sp12_h_r_14')
// (11, 13, 'sp4_h_r_19')
// (11, 15, 'sp4_h_r_28')
// (11, 17, 'sp4_r_v_b_42')
// (11, 18, 'sp4_r_v_b_31')
// (11, 19, 'sp4_r_v_b_18')
// (11, 20, 'sp4_h_r_36')
// (11, 20, 'sp4_r_v_b_7')
// (11, 21, 'sp4_r_v_b_42')
// (11, 22, 'local_g0_7')
// (11, 22, 'lutff_2/in_3')
// (11, 22, 'sp4_r_v_b_31')
// (11, 23, 'sp4_r_v_b_18')
// (11, 24, 'sp4_r_v_b_7')
// (12, 13, 'local_g2_6')
// (12, 13, 'lutff_2/in_0')
// (12, 13, 'sp12_h_r_17')
// (12, 13, 'sp4_h_r_30')
// (12, 15, 'sp4_h_r_41')
// (12, 16, 'sp4_r_v_b_41')
// (12, 16, 'sp4_v_t_42')
// (12, 17, 'sp4_r_v_b_28')
// (12, 17, 'sp4_v_b_42')
// (12, 18, 'sp4_r_v_b_17')
// (12, 18, 'sp4_v_b_31')
// (12, 19, 'local_g1_2')
// (12, 19, 'lutff_2/in_3')
// (12, 19, 'sp4_r_v_b_4')
// (12, 19, 'sp4_v_b_18')
// (12, 20, 'local_g0_7')
// (12, 20, 'lutff_2/in_3')
// (12, 20, 'sp4_h_l_36')
// (12, 20, 'sp4_h_r_7')
// (12, 20, 'sp4_v_b_7')
// (12, 20, 'sp4_v_t_42')
// (12, 21, 'sp4_v_b_42')
// (12, 22, 'sp4_v_b_31')
// (12, 23, 'sp4_v_b_18')
// (12, 24, 'sp4_v_b_7')
// (13, 13, 'sp12_h_r_18')
// (13, 13, 'sp4_h_r_43')
// (13, 14, 'sp4_r_v_b_46')
// (13, 15, 'sp4_h_l_41')
// (13, 15, 'sp4_h_r_4')
// (13, 15, 'sp4_r_v_b_35')
// (13, 15, 'sp4_v_t_41')
// (13, 16, 'local_g2_1')
// (13, 16, 'lutff_0/in_3')
// (13, 16, 'sp4_r_v_b_22')
// (13, 16, 'sp4_v_b_41')
// (13, 17, 'sp4_r_v_b_11')
// (13, 17, 'sp4_v_b_28')
// (13, 18, 'sp4_r_v_b_39')
// (13, 18, 'sp4_v_b_17')
// (13, 19, 'sp4_r_v_b_26')
// (13, 19, 'sp4_v_b_4')
// (13, 20, 'sp4_h_r_18')
// (13, 20, 'sp4_r_v_b_15')
// (13, 21, 'sp4_r_v_b_2')
// (14, 13, 'local_g0_5')
// (14, 13, 'lutff_2/in_3')
// (14, 13, 'sp12_h_r_21')
// (14, 13, 'sp4_h_l_43')
// (14, 13, 'sp4_v_t_46')
// (14, 14, 'sp4_v_b_46')
// (14, 15, 'sp4_h_r_17')
// (14, 15, 'sp4_v_b_35')
// (14, 16, 'sp4_v_b_22')
// (14, 17, 'sp4_v_b_11')
// (14, 17, 'sp4_v_t_39')
// (14, 18, 'sp4_v_b_39')
// (14, 19, 'sp4_v_b_26')
// (14, 20, 'sp4_h_r_31')
// (14, 20, 'sp4_v_b_15')
// (14, 21, 'local_g1_2')
// (14, 21, 'lutff_6/in_3')
// (14, 21, 'sp4_v_b_2')
// (15, 13, 'sp12_h_r_22')
// (15, 15, 'local_g3_4')
// (15, 15, 'lutff_2/in_3')
// (15, 15, 'sp4_h_r_28')
// (15, 17, 'local_g3_2')
// (15, 17, 'lutff_2/in_3')
// (15, 17, 'sp4_r_v_b_42')
// (15, 18, 'local_g0_7')
// (15, 18, 'lutff_2/in_3')
// (15, 18, 'sp4_r_v_b_31')
// (15, 19, 'sp4_r_v_b_18')
// (15, 19, 'sp4_r_v_b_40')
// (15, 20, 'sp4_h_r_42')
// (15, 20, 'sp4_r_v_b_29')
// (15, 20, 'sp4_r_v_b_7')
// (15, 21, 'sp4_r_v_b_16')
// (15, 22, 'sp4_r_v_b_5')
// (15, 23, 'sp4_r_v_b_36')
// (15, 24, 'sp4_r_v_b_25')
// (15, 25, 'sp4_r_v_b_12')
// (15, 26, 'sp4_r_v_b_1')
// (16, 1, 'sp12_v_t_22')
// (16, 2, 'sp12_v_b_22')
// (16, 3, 'sp12_v_b_21')
// (16, 4, 'sp12_v_b_18')
// (16, 5, 'sp12_v_b_17')
// (16, 6, 'sp12_v_b_14')
// (16, 7, 'sp12_v_b_13')
// (16, 8, 'sp12_v_b_10')
// (16, 9, 'sp12_v_b_9')
// (16, 10, 'sp12_v_b_6')
// (16, 11, 'local_g2_5')
// (16, 11, 'lutff_2/in_3')
// (16, 11, 'sp12_v_b_5')
// (16, 12, 'sp12_v_b_2')
// (16, 13, 'local_g1_1')
// (16, 13, 'lutff_1/in_1')
// (16, 13, 'sp12_h_l_22')
// (16, 13, 'sp12_h_r_1')
// (16, 13, 'sp12_v_b_1')
// (16, 13, 'sp12_v_t_22')
// (16, 14, 'sp12_v_b_22')
// (16, 15, 'sp12_v_b_21')
// (16, 15, 'sp4_h_r_41')
// (16, 16, 'local_g3_2')
// (16, 16, 'lutff_2/in_3')
// (16, 16, 'sp12_v_b_18')
// (16, 16, 'sp4_h_r_0')
// (16, 16, 'sp4_v_t_42')
// (16, 17, 'local_g2_1')
// (16, 17, 'lutff_2/in_3')
// (16, 17, 'sp12_v_b_17')
// (16, 17, 'sp4_v_b_42')
// (16, 18, 'local_g3_6')
// (16, 18, 'lutff_2/in_3')
// (16, 18, 'sp12_v_b_14')
// (16, 18, 'sp4_h_r_5')
// (16, 18, 'sp4_v_b_31')
// (16, 18, 'sp4_v_t_40')
// (16, 19, 'local_g2_5')
// (16, 19, 'lutff_0/in_3')
// (16, 19, 'sp12_v_b_13')
// (16, 19, 'sp4_v_b_18')
// (16, 19, 'sp4_v_b_40')
// (16, 20, 'sp12_v_b_10')
// (16, 20, 'sp4_h_l_42')
// (16, 20, 'sp4_h_r_7')
// (16, 20, 'sp4_v_b_29')
// (16, 20, 'sp4_v_b_7')
// (16, 21, 'local_g2_1')
// (16, 21, 'lutff_0/in_3')
// (16, 21, 'sp12_v_b_9')
// (16, 21, 'sp4_v_b_16')
// (16, 22, 'sp12_v_b_6')
// (16, 22, 'sp4_v_b_5')
// (16, 22, 'sp4_v_t_36')
// (16, 23, 'sp12_v_b_5')
// (16, 23, 'sp4_v_b_36')
// (16, 24, 'sp12_v_b_2')
// (16, 24, 'sp4_v_b_25')
// (16, 25, 'sp12_h_r_1')
// (16, 25, 'sp12_v_b_1')
// (16, 25, 'sp4_v_b_12')
// (16, 26, 'local_g1_1')
// (16, 26, 'lutff_5/in_3')
// (16, 26, 'sp4_v_b_1')
// (17, 10, 'sp4_r_v_b_39')
// (17, 11, 'sp4_r_v_b_26')
// (17, 12, 'sp4_r_v_b_15')
// (17, 13, 'sp12_h_r_2')
// (17, 13, 'sp4_r_v_b_2')
// (17, 15, 'sp4_h_l_41')
// (17, 16, 'sp4_h_r_13')
// (17, 18, 'sp4_h_r_16')
// (17, 20, 'sp4_h_r_18')
// (17, 25, 'sp12_h_r_2')
// (18, 9, 'sp4_v_t_39')
// (18, 10, 'sp4_v_b_39')
// (18, 11, 'local_g3_2')
// (18, 11, 'lutff_2/in_3')
// (18, 11, 'sp4_v_b_26')
// (18, 12, 'local_g0_7')
// (18, 12, 'lutff_2/in_3')
// (18, 12, 'sp4_v_b_15')
// (18, 13, 'sp12_h_r_5')
// (18, 13, 'sp4_h_r_2')
// (18, 13, 'sp4_v_b_2')
// (18, 16, 'sp4_h_r_24')
// (18, 18, 'sp4_h_r_29')
// (18, 20, 'sp4_h_r_31')
// (18, 25, 'sp12_h_r_5')
// (19, 10, 'local_g3_1')
// (19, 10, 'lutff_2/in_0')
// (19, 10, 'sp4_r_v_b_41')
// (19, 11, 'local_g1_4')
// (19, 11, 'lutff_2/in_3')
// (19, 11, 'sp4_r_v_b_28')
// (19, 12, 'sp4_r_v_b_17')
// (19, 13, 'sp12_h_r_6')
// (19, 13, 'sp4_h_r_15')
// (19, 13, 'sp4_r_v_b_4')
// (19, 16, 'local_g2_5')
// (19, 16, 'lutff_2/in_3')
// (19, 16, 'sp4_h_r_37')
// (19, 17, 'sp4_r_v_b_36')
// (19, 18, 'sp4_h_r_40')
// (19, 18, 'sp4_r_v_b_25')
// (19, 19, 'local_g2_4')
// (19, 19, 'lutff_1/in_3')
// (19, 19, 'sp4_r_v_b_12')
// (19, 20, 'sp4_h_r_42')
// (19, 20, 'sp4_r_v_b_1')
// (19, 21, 'sp4_r_v_b_37')
// (19, 22, 'sp4_r_v_b_24')
// (19, 23, 'sp4_r_v_b_13')
// (19, 24, 'sp4_r_v_b_0')
// (19, 25, 'local_g1_6')
// (19, 25, 'lutff_2/in_3')
// (19, 25, 'sp12_h_r_6')
// (20, 9, 'sp4_v_t_41')
// (20, 10, 'sp4_v_b_41')
// (20, 11, 'local_g2_4')
// (20, 11, 'lutff_1/in_3')
// (20, 11, 'sp4_v_b_28')
// (20, 12, 'local_g0_1')
// (20, 12, 'lutff_2/in_1')
// (20, 12, 'sp4_v_b_17')
// (20, 13, 'local_g3_2')
// (20, 13, 'lutff_7/in_0')
// (20, 13, 'sp12_h_r_9')
// (20, 13, 'sp4_h_r_26')
// (20, 13, 'sp4_h_r_4')
// (20, 13, 'sp4_v_b_4')
// (20, 16, 'local_g0_3')
// (20, 16, 'lutff_2/in_3')
// (20, 16, 'sp4_h_l_37')
// (20, 16, 'sp4_h_r_3')
// (20, 16, 'sp4_v_t_36')
// (20, 17, 'local_g2_4')
// (20, 17, 'lutff_5/in_3')
// (20, 17, 'sp4_v_b_36')
// (20, 18, 'local_g3_1')
// (20, 18, 'lutff_6/in_0')
// (20, 18, 'sp4_h_l_40')
// (20, 18, 'sp4_h_r_8')
// (20, 18, 'sp4_v_b_25')
// (20, 19, 'local_g1_4')
// (20, 19, 'lutff_2/in_3')
// (20, 19, 'sp4_v_b_12')
// (20, 20, 'local_g0_1')
// (20, 20, 'lutff_2/in_1')
// (20, 20, 'sp4_h_l_42')
// (20, 20, 'sp4_h_r_10')
// (20, 20, 'sp4_v_b_1')
// (20, 20, 'sp4_v_t_37')
// (20, 21, 'sp4_v_b_37')
// (20, 22, 'sp4_v_b_24')
// (20, 23, 'local_g1_5')
// (20, 23, 'lutff_5/in_3')
// (20, 23, 'sp4_v_b_13')
// (20, 24, 'sp4_v_b_0')
// (20, 25, 'local_g0_1')
// (20, 25, 'lutff_2/in_1')
// (20, 25, 'sp12_h_r_9')
// (21, 10, 'sp4_r_v_b_39')
// (21, 11, 'local_g0_2')
// (21, 11, 'lutff_2/in_0')
// (21, 11, 'sp4_r_v_b_26')
// (21, 12, 'local_g2_7')
// (21, 12, 'lutff_2/in_3')
// (21, 12, 'sp4_r_v_b_15')
// (21, 13, 'sp12_h_r_10')
// (21, 13, 'sp4_h_r_17')
// (21, 13, 'sp4_h_r_39')
// (21, 13, 'sp4_r_v_b_2')
// (21, 14, 'sp4_r_v_b_43')
// (21, 15, 'sp4_r_v_b_30')
// (21, 16, 'local_g0_6')
// (21, 16, 'lutff_0/in_0')
// (21, 16, 'sp4_h_r_14')
// (21, 16, 'sp4_r_v_b_19')
// (21, 17, 'sp4_r_v_b_6')
// (21, 18, 'local_g0_5')
// (21, 18, 'lutff_2/in_3')
// (21, 18, 'sp4_h_r_21')
// (21, 20, 'local_g0_7')
// (21, 20, 'lutff_2/in_3')
// (21, 20, 'sp4_h_r_23')
// (21, 22, 'sp4_r_v_b_46')
// (21, 23, 'sp4_r_v_b_35')
// (21, 24, 'sp4_r_v_b_22')
// (21, 25, 'sp12_h_r_10')
// (21, 25, 'sp4_r_v_b_11')
// (22, 9, 'sp4_v_t_39')
// (22, 10, 'sp4_v_b_39')
// (22, 11, 'sp4_v_b_26')
// (22, 12, 'local_g0_7')
// (22, 12, 'lutff_2/in_3')
// (22, 12, 'sp4_v_b_15')
// (22, 13, 'sp12_h_r_13')
// (22, 13, 'sp4_h_l_39')
// (22, 13, 'sp4_h_r_28')
// (22, 13, 'sp4_h_r_6')
// (22, 13, 'sp4_v_b_2')
// (22, 13, 'sp4_v_t_43')
// (22, 14, 'local_g2_3')
// (22, 14, 'lutff_2/in_3')
// (22, 14, 'sp4_v_b_43')
// (22, 15, 'sp4_v_b_30')
// (22, 16, 'sp4_h_r_27')
// (22, 16, 'sp4_v_b_19')
// (22, 17, 'sp4_v_b_6')
// (22, 18, 'sp4_h_r_32')
// (22, 20, 'local_g3_2')
// (22, 20, 'lutff_5/in_0')
// (22, 20, 'sp4_h_r_34')
// (22, 21, 'local_g1_4')
// (22, 21, 'lutff_2/in_3')
// (22, 21, 'sp4_h_r_4')
// (22, 21, 'sp4_v_t_46')
// (22, 22, 'sp4_v_b_46')
// (22, 23, 'local_g2_3')
// (22, 23, 'lutff_2/in_3')
// (22, 23, 'sp4_v_b_35')
// (22, 24, 'sp4_v_b_22')
// (22, 25, 'sp12_h_r_13')
// (22, 25, 'sp4_h_r_6')
// (22, 25, 'sp4_v_b_11')
// (23, 10, 'sp4_r_v_b_41')
// (23, 11, 'sp4_r_v_b_28')
// (23, 12, 'local_g3_1')
// (23, 12, 'lutff_2/in_0')
// (23, 12, 'sp4_r_v_b_17')
// (23, 13, 'sp12_h_r_14')
// (23, 13, 'sp4_h_r_19')
// (23, 13, 'sp4_h_r_41')
// (23, 13, 'sp4_r_v_b_4')
// (23, 14, 'local_g3_1')
// (23, 14, 'lutff_2/in_0')
// (23, 14, 'sp4_r_v_b_41')
// (23, 14, 'sp4_r_v_b_44')
// (23, 15, 'local_g2_1')
// (23, 15, 'lutff_2/in_3')
// (23, 15, 'sp4_r_v_b_28')
// (23, 15, 'sp4_r_v_b_33')
// (23, 16, 'local_g3_4')
// (23, 16, 'lutff_2/in_3')
// (23, 16, 'sp4_h_r_38')
// (23, 16, 'sp4_r_v_b_17')
// (23, 16, 'sp4_r_v_b_20')
// (23, 17, 'sp4_r_v_b_4')
// (23, 17, 'sp4_r_v_b_9')
// (23, 18, 'sp4_h_r_45')
// (23, 20, 'local_g2_7')
// (23, 20, 'lutff_2/in_3')
// (23, 20, 'sp4_h_r_47')
// (23, 21, 'sp4_h_r_17')
// (23, 25, 'sp12_h_r_14')
// (23, 25, 'sp4_h_r_19')
// (24, 9, 'sp4_v_t_41')
// (24, 10, 'sp4_v_b_41')
// (24, 11, 'sp4_v_b_28')
// (24, 12, 'sp4_v_b_17')
// (24, 13, 'local_g0_1')
// (24, 13, 'lutff_0/in_1')
// (24, 13, 'sp12_h_r_17')
// (24, 13, 'sp4_h_l_41')
// (24, 13, 'sp4_h_r_30')
// (24, 13, 'sp4_v_b_4')
// (24, 13, 'sp4_v_t_41')
// (24, 13, 'sp4_v_t_44')
// (24, 14, 'local_g3_4')
// (24, 14, 'lutff_2/in_3')
// (24, 14, 'sp4_v_b_41')
// (24, 14, 'sp4_v_b_44')
// (24, 15, 'sp4_v_b_28')
// (24, 15, 'sp4_v_b_33')
// (24, 16, 'local_g1_4')
// (24, 16, 'lutff_0/in_3')
// (24, 16, 'sp4_h_l_38')
// (24, 16, 'sp4_v_b_17')
// (24, 16, 'sp4_v_b_20')
// (24, 17, 'local_g1_4')
// (24, 17, 'lutff_2/in_3')
// (24, 17, 'sp4_v_b_4')
// (24, 17, 'sp4_v_b_9')
// (24, 18, 'sp4_h_l_45')
// (24, 20, 'sp4_h_l_47')
// (24, 21, 'sp4_h_r_28')
// (24, 25, 'sp12_h_r_17')
// (24, 25, 'sp4_h_r_30')
// (25, 13, 'sp12_h_r_18')
// (25, 13, 'sp4_h_r_43')
// (25, 21, 'sp4_h_r_41')
// (25, 25, 'sp12_h_r_18')
// (25, 25, 'sp4_h_r_43')
// (26, 13, 'sp12_h_r_21')
// (26, 13, 'sp4_h_l_43')
// (26, 21, 'sp4_h_l_41')
// (26, 25, 'sp12_h_r_21')
// (26, 25, 'sp4_h_l_43')
// (27, 13, 'sp12_h_r_22')
// (27, 25, 'sp12_h_r_22')
// (28, 13, 'sp12_h_l_22')
// (28, 25, 'sp12_h_l_22')

reg n45 = 0;
// (4, 16, 'neigh_op_tnr_0')
// (4, 17, 'neigh_op_rgt_0')
// (4, 18, 'neigh_op_bnr_0')
// (5, 13, 'sp12_v_t_23')
// (5, 14, 'sp12_v_b_23')
// (5, 15, 'sp12_v_b_20')
// (5, 16, 'neigh_op_top_0')
// (5, 16, 'sp12_v_b_19')
// (5, 17, 'local_g3_0')
// (5, 17, 'lutff_0/in_1')
// (5, 17, 'lutff_0/out')
// (5, 17, 'sp12_v_b_16')
// (5, 18, 'neigh_op_bot_0')
// (5, 18, 'sp12_v_b_15')
// (5, 19, 'sp12_v_b_12')
// (5, 20, 'sp12_v_b_11')
// (5, 21, 'sp12_v_b_8')
// (5, 22, 'sp12_v_b_7')
// (5, 23, 'sp12_v_b_4')
// (5, 24, 'sp12_v_b_3')
// (5, 25, 'sp12_h_r_0')
// (5, 25, 'sp12_v_b_0')
// (6, 16, 'neigh_op_tnl_0')
// (6, 17, 'neigh_op_lft_0')
// (6, 18, 'neigh_op_bnl_0')
// (6, 25, 'sp12_h_r_3')
// (7, 25, 'sp12_h_r_4')
// (8, 25, 'sp12_h_r_7')
// (9, 25, 'sp12_h_r_8')
// (10, 25, 'sp12_h_r_11')
// (11, 25, 'sp12_h_r_12')
// (12, 25, 'sp12_h_r_15')
// (13, 25, 'sp12_h_r_16')
// (14, 25, 'sp12_h_r_19')
// (15, 25, 'sp12_h_r_20')
// (16, 24, 'sp4_r_v_b_47')
// (16, 25, 'sp12_h_r_23')
// (16, 25, 'sp4_r_v_b_34')
// (16, 26, 'sp4_r_v_b_23')
// (16, 27, 'sp4_r_v_b_10')
// (17, 23, 'sp4_h_r_10')
// (17, 23, 'sp4_v_t_47')
// (17, 24, 'sp4_v_b_47')
// (17, 25, 'sp12_h_l_23')
// (17, 25, 'sp12_v_t_23')
// (17, 25, 'sp4_v_b_34')
// (17, 26, 'sp12_v_b_23')
// (17, 26, 'sp4_v_b_23')
// (17, 27, 'sp12_v_b_20')
// (17, 27, 'sp4_v_b_10')
// (17, 28, 'sp12_v_b_19')
// (17, 29, 'sp12_v_b_16')
// (17, 30, 'sp12_v_b_15')
// (17, 31, 'sp12_v_b_12')
// (17, 32, 'sp12_v_b_11')
// (17, 33, 'span12_vert_8')
// (18, 23, 'local_g1_7')
// (18, 23, 'lutff_0/in_0')
// (18, 23, 'sp4_h_r_23')
// (19, 23, 'sp4_h_r_34')
// (20, 23, 'sp4_h_r_47')
// (21, 23, 'sp4_h_l_47')

reg n46 = 0;
// (4, 16, 'neigh_op_tnr_1')
// (4, 17, 'neigh_op_rgt_1')
// (4, 18, 'neigh_op_bnr_1')
// (5, 16, 'neigh_op_top_1')
// (5, 17, 'local_g3_1')
// (5, 17, 'lutff_1/in_1')
// (5, 17, 'lutff_1/out')
// (5, 17, 'sp4_h_r_2')
// (5, 18, 'neigh_op_bot_1')
// (6, 16, 'neigh_op_tnl_1')
// (6, 17, 'neigh_op_lft_1')
// (6, 17, 'sp4_h_r_15')
// (6, 18, 'neigh_op_bnl_1')
// (7, 17, 'sp4_h_r_26')
// (8, 17, 'sp4_h_r_39')
// (8, 18, 'sp4_r_v_b_42')
// (8, 19, 'sp4_r_v_b_31')
// (8, 20, 'sp4_r_v_b_18')
// (8, 21, 'sp4_r_v_b_7')
// (9, 17, 'sp4_h_l_39')
// (9, 17, 'sp4_v_t_42')
// (9, 18, 'sp4_v_b_42')
// (9, 19, 'sp4_v_b_31')
// (9, 20, 'sp4_v_b_18')
// (9, 21, 'sp4_h_r_1')
// (9, 21, 'sp4_v_b_7')
// (10, 21, 'sp4_h_r_12')
// (11, 21, 'sp4_h_r_25')
// (12, 21, 'sp4_h_r_36')
// (13, 21, 'sp4_h_l_36')
// (13, 21, 'sp4_h_r_1')
// (14, 21, 'sp4_h_r_12')
// (15, 21, 'sp4_h_r_25')
// (16, 21, 'sp4_h_r_36')
// (17, 21, 'sp4_h_l_36')
// (17, 21, 'sp4_h_r_4')
// (18, 21, 'local_g1_1')
// (18, 21, 'lutff_7/in_1')
// (18, 21, 'sp4_h_r_17')
// (19, 21, 'sp4_h_r_28')
// (20, 21, 'sp4_h_r_41')
// (21, 21, 'sp4_h_l_41')

reg n47 = 0;
// (4, 16, 'neigh_op_tnr_3')
// (4, 17, 'neigh_op_rgt_3')
// (4, 18, 'neigh_op_bnr_3')
// (5, 16, 'neigh_op_top_3')
// (5, 16, 'sp12_v_t_22')
// (5, 17, 'local_g1_3')
// (5, 17, 'lutff_3/in_1')
// (5, 17, 'lutff_3/out')
// (5, 17, 'sp12_v_b_22')
// (5, 18, 'neigh_op_bot_3')
// (5, 18, 'sp12_v_b_21')
// (5, 19, 'sp12_v_b_18')
// (5, 20, 'sp12_v_b_17')
// (5, 21, 'sp12_v_b_14')
// (5, 22, 'sp12_v_b_13')
// (5, 23, 'sp12_v_b_10')
// (5, 24, 'sp12_v_b_9')
// (5, 25, 'sp12_v_b_6')
// (5, 26, 'sp12_v_b_5')
// (5, 27, 'sp12_v_b_2')
// (5, 28, 'sp12_h_r_1')
// (5, 28, 'sp12_v_b_1')
// (6, 16, 'neigh_op_tnl_3')
// (6, 17, 'neigh_op_lft_3')
// (6, 18, 'neigh_op_bnl_3')
// (6, 28, 'sp12_h_r_2')
// (7, 28, 'sp12_h_r_5')
// (8, 28, 'sp12_h_r_6')
// (9, 28, 'sp12_h_r_9')
// (10, 28, 'sp12_h_r_10')
// (11, 28, 'sp12_h_r_13')
// (12, 28, 'sp12_h_r_14')
// (13, 28, 'sp12_h_r_17')
// (14, 28, 'sp12_h_r_18')
// (15, 28, 'sp12_h_r_21')
// (15, 28, 'sp4_h_r_10')
// (16, 28, 'sp12_h_r_22')
// (16, 28, 'sp4_h_r_23')
// (17, 28, 'sp12_h_l_22')
// (17, 28, 'sp4_h_r_34')
// (18, 21, 'sp4_r_v_b_36')
// (18, 22, 'sp4_r_v_b_25')
// (18, 23, 'local_g2_4')
// (18, 23, 'lutff_5/in_3')
// (18, 23, 'sp4_r_v_b_12')
// (18, 24, 'sp4_r_v_b_1')
// (18, 25, 'sp4_r_v_b_47')
// (18, 26, 'sp4_r_v_b_34')
// (18, 27, 'sp4_r_v_b_23')
// (18, 28, 'sp4_h_r_47')
// (18, 28, 'sp4_r_v_b_10')
// (19, 20, 'sp4_v_t_36')
// (19, 21, 'sp4_v_b_36')
// (19, 22, 'sp4_v_b_25')
// (19, 23, 'sp4_v_b_12')
// (19, 24, 'sp4_v_b_1')
// (19, 24, 'sp4_v_t_47')
// (19, 25, 'sp4_v_b_47')
// (19, 26, 'sp4_v_b_34')
// (19, 27, 'sp4_v_b_23')
// (19, 28, 'sp4_h_l_47')
// (19, 28, 'sp4_v_b_10')

reg n48 = 0;
// (4, 16, 'neigh_op_tnr_4')
// (4, 17, 'neigh_op_rgt_4')
// (4, 18, 'neigh_op_bnr_4')
// (5, 16, 'neigh_op_top_4')
// (5, 17, 'local_g3_4')
// (5, 17, 'lutff_4/in_1')
// (5, 17, 'lutff_4/out')
// (5, 17, 'sp4_h_r_8')
// (5, 18, 'neigh_op_bot_4')
// (6, 16, 'neigh_op_tnl_4')
// (6, 17, 'neigh_op_lft_4')
// (6, 17, 'sp4_h_r_21')
// (6, 18, 'neigh_op_bnl_4')
// (7, 17, 'sp4_h_r_32')
// (8, 17, 'sp4_h_r_45')
// (9, 17, 'sp4_h_l_45')
// (9, 17, 'sp4_h_r_4')
// (10, 17, 'sp4_h_r_17')
// (11, 17, 'sp4_h_r_28')
// (12, 17, 'sp4_h_r_41')
// (12, 18, 'sp4_r_v_b_44')
// (12, 19, 'sp4_r_v_b_33')
// (12, 20, 'sp4_r_v_b_20')
// (12, 21, 'sp4_r_v_b_9')
// (13, 17, 'sp4_h_l_41')
// (13, 17, 'sp4_v_t_44')
// (13, 18, 'sp4_v_b_44')
// (13, 19, 'sp4_v_b_33')
// (13, 20, 'sp4_v_b_20')
// (13, 21, 'sp4_h_r_9')
// (13, 21, 'sp4_v_b_9')
// (14, 21, 'sp4_h_r_20')
// (15, 21, 'sp4_h_r_33')
// (16, 21, 'sp4_h_r_44')
// (17, 21, 'sp4_h_l_44')
// (17, 21, 'sp4_h_r_9')
// (18, 21, 'local_g0_4')
// (18, 21, 'lutff_5/in_1')
// (18, 21, 'sp4_h_r_20')
// (19, 21, 'sp4_h_r_33')
// (20, 21, 'sp4_h_r_44')
// (21, 21, 'sp4_h_l_44')

reg n49 = 0;
// (4, 16, 'neigh_op_tnr_5')
// (4, 17, 'neigh_op_rgt_5')
// (4, 18, 'neigh_op_bnr_5')
// (5, 16, 'neigh_op_top_5')
// (5, 16, 'sp4_r_v_b_38')
// (5, 17, 'local_g1_5')
// (5, 17, 'lutff_5/in_1')
// (5, 17, 'lutff_5/out')
// (5, 17, 'sp4_r_v_b_27')
// (5, 18, 'neigh_op_bot_5')
// (5, 18, 'sp4_r_v_b_14')
// (5, 19, 'sp4_r_v_b_3')
// (6, 15, 'sp4_v_t_38')
// (6, 16, 'neigh_op_tnl_5')
// (6, 16, 'sp4_v_b_38')
// (6, 17, 'neigh_op_lft_5')
// (6, 17, 'sp4_v_b_27')
// (6, 18, 'neigh_op_bnl_5')
// (6, 18, 'sp4_v_b_14')
// (6, 19, 'sp4_h_r_9')
// (6, 19, 'sp4_v_b_3')
// (7, 19, 'sp4_h_r_20')
// (8, 19, 'sp4_h_r_33')
// (9, 19, 'sp4_h_r_44')
// (10, 19, 'sp4_h_l_44')
// (10, 19, 'sp4_h_r_9')
// (11, 19, 'sp4_h_r_20')
// (12, 19, 'sp4_h_r_33')
// (13, 19, 'sp4_h_r_44')
// (14, 19, 'sp4_h_l_44')
// (14, 19, 'sp4_h_r_5')
// (15, 19, 'sp4_h_r_16')
// (16, 19, 'sp4_h_r_29')
// (17, 19, 'sp4_h_r_40')
// (17, 20, 'sp4_r_v_b_47')
// (17, 21, 'sp4_r_v_b_34')
// (17, 22, 'sp4_r_v_b_23')
// (17, 23, 'sp4_r_v_b_10')
// (18, 19, 'sp4_h_l_40')
// (18, 19, 'sp4_v_t_47')
// (18, 20, 'sp4_v_b_47')
// (18, 21, 'sp4_v_b_34')
// (18, 22, 'sp4_v_b_23')
// (18, 23, 'local_g1_2')
// (18, 23, 'lutff_4/in_3')
// (18, 23, 'sp4_v_b_10')

reg n50 = 0;
// (4, 16, 'neigh_op_tnr_6')
// (4, 17, 'neigh_op_rgt_6')
// (4, 18, 'neigh_op_bnr_6')
// (5, 11, 'sp12_v_t_23')
// (5, 12, 'sp12_v_b_23')
// (5, 13, 'sp12_v_b_20')
// (5, 14, 'sp12_v_b_19')
// (5, 15, 'sp12_v_b_16')
// (5, 16, 'neigh_op_top_6')
// (5, 16, 'sp12_v_b_15')
// (5, 17, 'local_g1_6')
// (5, 17, 'lutff_6/in_1')
// (5, 17, 'lutff_6/out')
// (5, 17, 'sp12_v_b_12')
// (5, 18, 'neigh_op_bot_6')
// (5, 18, 'sp12_v_b_11')
// (5, 19, 'sp12_v_b_8')
// (5, 20, 'sp12_v_b_7')
// (5, 21, 'sp12_v_b_4')
// (5, 22, 'sp12_v_b_3')
// (5, 23, 'sp12_h_r_0')
// (5, 23, 'sp12_v_b_0')
// (6, 16, 'neigh_op_tnl_6')
// (6, 17, 'neigh_op_lft_6')
// (6, 18, 'neigh_op_bnl_6')
// (6, 23, 'sp12_h_r_3')
// (7, 23, 'sp12_h_r_4')
// (8, 23, 'sp12_h_r_7')
// (9, 23, 'sp12_h_r_8')
// (10, 23, 'sp12_h_r_11')
// (11, 23, 'sp12_h_r_12')
// (12, 23, 'sp12_h_r_15')
// (13, 23, 'sp12_h_r_16')
// (14, 23, 'sp12_h_r_19')
// (15, 23, 'sp12_h_r_20')
// (16, 23, 'sp12_h_r_23')
// (17, 23, 'sp12_h_l_23')
// (17, 23, 'sp12_h_r_0')
// (18, 23, 'local_g1_3')
// (18, 23, 'lutff_1/in_3')
// (18, 23, 'sp12_h_r_3')
// (19, 23, 'sp12_h_r_4')
// (20, 23, 'sp12_h_r_7')
// (21, 23, 'sp12_h_r_8')
// (22, 23, 'sp12_h_r_11')
// (23, 23, 'sp12_h_r_12')
// (24, 23, 'sp12_h_r_15')
// (25, 23, 'sp12_h_r_16')
// (26, 23, 'sp12_h_r_19')
// (27, 23, 'sp12_h_r_20')
// (28, 23, 'sp12_h_r_23')
// (29, 23, 'sp12_h_l_23')

reg n51 = 0;
// (4, 16, 'sp12_h_r_1')
// (5, 16, 'sp12_h_r_2')
// (6, 15, 'neigh_op_tnr_7')
// (6, 16, 'neigh_op_rgt_7')
// (6, 16, 'sp12_h_r_5')
// (6, 17, 'neigh_op_bnr_7')
// (7, 15, 'neigh_op_top_7')
// (7, 16, 'lutff_7/out')
// (7, 16, 'sp12_h_r_6')
// (7, 17, 'neigh_op_bot_7')
// (8, 15, 'neigh_op_tnl_7')
// (8, 16, 'neigh_op_lft_7')
// (8, 16, 'sp12_h_r_9')
// (8, 17, 'neigh_op_bnl_7')
// (9, 16, 'sp12_h_r_10')
// (10, 16, 'sp12_h_r_13')
// (11, 16, 'local_g0_6')
// (11, 16, 'lutff_4/in_0')
// (11, 16, 'lutff_5/in_3')
// (11, 16, 'lutff_7/in_3')
// (11, 16, 'sp12_h_r_14')
// (12, 16, 'sp12_h_r_17')
// (13, 16, 'sp12_h_r_18')
// (14, 16, 'sp12_h_r_21')
// (15, 16, 'sp12_h_r_22')
// (16, 16, 'sp12_h_l_22')

reg n52 = 0;
// (4, 17, 'neigh_op_tnr_0')
// (4, 18, 'neigh_op_rgt_0')
// (4, 18, 'sp4_h_r_5')
// (4, 19, 'neigh_op_bnr_0')
// (5, 17, 'neigh_op_top_0')
// (5, 18, 'local_g3_0')
// (5, 18, 'lutff_0/in_1')
// (5, 18, 'lutff_0/out')
// (5, 18, 'sp4_h_r_16')
// (5, 19, 'neigh_op_bot_0')
// (6, 17, 'neigh_op_tnl_0')
// (6, 18, 'neigh_op_lft_0')
// (6, 18, 'sp4_h_r_29')
// (6, 19, 'neigh_op_bnl_0')
// (7, 18, 'sp4_h_r_40')
// (8, 18, 'sp4_h_l_40')
// (8, 18, 'sp4_h_r_5')
// (9, 18, 'sp4_h_r_16')
// (10, 18, 'sp4_h_r_29')
// (11, 18, 'sp4_h_r_40')
// (12, 18, 'sp4_h_l_40')
// (12, 18, 'sp4_h_r_1')
// (13, 18, 'sp4_h_r_12')
// (14, 18, 'sp4_h_r_25')
// (15, 18, 'sp4_h_r_36')
// (15, 19, 'sp4_r_v_b_36')
// (15, 20, 'sp4_r_v_b_25')
// (15, 21, 'sp4_r_v_b_12')
// (15, 22, 'sp4_r_v_b_1')
// (16, 18, 'sp4_h_l_36')
// (16, 18, 'sp4_v_t_36')
// (16, 19, 'sp4_v_b_36')
// (16, 20, 'sp4_v_b_25')
// (16, 21, 'sp4_v_b_12')
// (16, 22, 'local_g0_1')
// (16, 22, 'lutff_1/in_2')
// (16, 22, 'sp4_v_b_1')

reg n53 = 0;
// (4, 17, 'neigh_op_tnr_1')
// (4, 18, 'neigh_op_rgt_1')
// (4, 19, 'neigh_op_bnr_1')
// (5, 17, 'neigh_op_top_1')
// (5, 18, 'local_g3_1')
// (5, 18, 'lutff_1/in_1')
// (5, 18, 'lutff_1/out')
// (5, 18, 'sp4_h_r_2')
// (5, 19, 'neigh_op_bot_1')
// (6, 17, 'neigh_op_tnl_1')
// (6, 18, 'neigh_op_lft_1')
// (6, 18, 'sp4_h_r_15')
// (6, 19, 'neigh_op_bnl_1')
// (7, 18, 'sp4_h_r_26')
// (8, 18, 'sp4_h_r_39')
// (8, 19, 'sp4_r_v_b_39')
// (8, 20, 'sp4_r_v_b_26')
// (8, 21, 'sp4_r_v_b_15')
// (8, 22, 'sp4_r_v_b_2')
// (9, 18, 'sp4_h_l_39')
// (9, 18, 'sp4_v_t_39')
// (9, 19, 'sp4_v_b_39')
// (9, 20, 'sp4_v_b_26')
// (9, 21, 'sp4_v_b_15')
// (9, 22, 'sp4_h_r_8')
// (9, 22, 'sp4_v_b_2')
// (10, 22, 'sp4_h_r_21')
// (11, 22, 'sp4_h_r_32')
// (12, 22, 'sp4_h_r_45')
// (13, 22, 'sp4_h_l_45')
// (13, 22, 'sp4_h_r_8')
// (14, 22, 'sp4_h_r_21')
// (15, 22, 'sp4_h_r_32')
// (16, 22, 'local_g2_5')
// (16, 22, 'lutff_2/in_1')
// (16, 22, 'sp4_h_r_45')
// (17, 22, 'sp4_h_l_45')

reg n54 = 0;
// (4, 17, 'neigh_op_tnr_2')
// (4, 18, 'neigh_op_rgt_2')
// (4, 19, 'neigh_op_bnr_2')
// (5, 17, 'neigh_op_top_2')
// (5, 18, 'local_g1_2')
// (5, 18, 'lutff_2/in_1')
// (5, 18, 'lutff_2/out')
// (5, 18, 'sp4_r_v_b_37')
// (5, 19, 'neigh_op_bot_2')
// (5, 19, 'sp4_r_v_b_24')
// (5, 20, 'sp4_r_v_b_13')
// (5, 21, 'sp4_r_v_b_0')
// (6, 17, 'neigh_op_tnl_2')
// (6, 17, 'sp4_v_t_37')
// (6, 18, 'neigh_op_lft_2')
// (6, 18, 'sp4_v_b_37')
// (6, 19, 'neigh_op_bnl_2')
// (6, 19, 'sp4_v_b_24')
// (6, 20, 'sp4_v_b_13')
// (6, 21, 'sp4_h_r_6')
// (6, 21, 'sp4_v_b_0')
// (7, 21, 'sp4_h_r_19')
// (8, 21, 'sp4_h_r_30')
// (9, 21, 'sp4_h_r_43')
// (10, 21, 'sp4_h_l_43')
// (10, 21, 'sp4_h_r_2')
// (11, 21, 'sp4_h_r_15')
// (12, 21, 'sp4_h_r_26')
// (13, 21, 'sp4_h_r_39')
// (14, 21, 'sp4_h_l_39')
// (14, 21, 'sp4_h_r_10')
// (15, 21, 'sp4_h_r_23')
// (16, 21, 'sp4_h_r_34')
// (17, 21, 'sp4_h_r_47')
// (17, 22, 'sp4_r_v_b_47')
// (17, 23, 'sp4_r_v_b_34')
// (17, 24, 'sp4_r_v_b_23')
// (17, 25, 'sp4_r_v_b_10')
// (18, 21, 'sp4_h_l_47')
// (18, 21, 'sp4_v_t_47')
// (18, 22, 'sp4_v_b_47')
// (18, 23, 'local_g2_2')
// (18, 23, 'lutff_2/in_0')
// (18, 23, 'sp4_v_b_34')
// (18, 24, 'sp4_v_b_23')
// (18, 25, 'sp4_v_b_10')

reg n55 = 0;
// (4, 17, 'neigh_op_tnr_3')
// (4, 18, 'neigh_op_rgt_3')
// (4, 19, 'neigh_op_bnr_3')
// (5, 16, 'sp4_r_v_b_47')
// (5, 17, 'neigh_op_top_3')
// (5, 17, 'sp4_r_v_b_34')
// (5, 18, 'local_g1_3')
// (5, 18, 'lutff_3/in_1')
// (5, 18, 'lutff_3/out')
// (5, 18, 'sp4_r_v_b_23')
// (5, 19, 'neigh_op_bot_3')
// (5, 19, 'sp4_r_v_b_10')
// (6, 15, 'sp4_v_t_47')
// (6, 16, 'sp4_v_b_47')
// (6, 17, 'neigh_op_tnl_3')
// (6, 17, 'sp4_v_b_34')
// (6, 18, 'neigh_op_lft_3')
// (6, 18, 'sp4_v_b_23')
// (6, 19, 'neigh_op_bnl_3')
// (6, 19, 'sp4_h_r_10')
// (6, 19, 'sp4_v_b_10')
// (7, 19, 'sp4_h_r_23')
// (8, 19, 'sp4_h_r_34')
// (9, 19, 'sp4_h_r_47')
// (10, 19, 'sp4_h_l_47')
// (10, 19, 'sp4_h_r_1')
// (11, 19, 'sp4_h_r_12')
// (12, 19, 'sp4_h_r_25')
// (13, 19, 'sp4_h_r_36')
// (14, 19, 'sp4_h_l_36')
// (14, 19, 'sp4_h_r_4')
// (15, 19, 'sp4_h_r_17')
// (16, 19, 'sp4_h_r_28')
// (17, 19, 'sp4_h_r_41')
// (17, 20, 'sp4_r_v_b_41')
// (17, 21, 'sp4_r_v_b_28')
// (17, 22, 'sp4_r_v_b_17')
// (17, 23, 'sp4_r_v_b_4')
// (18, 19, 'sp4_h_l_41')
// (18, 19, 'sp4_v_t_41')
// (18, 20, 'sp4_v_b_41')
// (18, 21, 'sp4_v_b_28')
// (18, 22, 'sp4_v_b_17')
// (18, 23, 'local_g0_4')
// (18, 23, 'lutff_3/in_1')
// (18, 23, 'sp4_v_b_4')

reg n56 = 0;
// (4, 17, 'neigh_op_tnr_4')
// (4, 18, 'neigh_op_rgt_4')
// (4, 19, 'neigh_op_bnr_4')
// (5, 17, 'neigh_op_top_4')
// (5, 18, 'local_g1_4')
// (5, 18, 'lutff_4/in_1')
// (5, 18, 'lutff_4/out')
// (5, 18, 'sp12_h_r_0')
// (5, 19, 'neigh_op_bot_4')
// (6, 17, 'neigh_op_tnl_4')
// (6, 18, 'neigh_op_lft_4')
// (6, 18, 'sp12_h_r_3')
// (6, 19, 'neigh_op_bnl_4')
// (7, 18, 'sp12_h_r_4')
// (8, 18, 'sp12_h_r_7')
// (9, 18, 'sp12_h_r_8')
// (10, 18, 'sp12_h_r_11')
// (11, 18, 'sp12_h_r_12')
// (12, 18, 'sp12_h_r_15')
// (13, 18, 'sp12_h_r_16')
// (14, 18, 'sp12_h_r_19')
// (14, 18, 'sp4_h_r_11')
// (15, 18, 'sp12_h_r_20')
// (15, 18, 'sp4_h_r_22')
// (16, 18, 'sp12_h_r_23')
// (16, 18, 'sp4_h_r_35')
// (17, 18, 'sp12_h_l_23')
// (17, 18, 'sp4_h_r_46')
// (17, 19, 'sp4_r_v_b_46')
// (17, 20, 'sp4_r_v_b_35')
// (17, 21, 'sp4_r_v_b_22')
// (17, 22, 'sp4_r_v_b_11')
// (18, 18, 'sp4_h_l_46')
// (18, 18, 'sp4_v_t_46')
// (18, 19, 'sp4_v_b_46')
// (18, 20, 'sp4_v_b_35')
// (18, 21, 'local_g0_6')
// (18, 21, 'lutff_6/in_0')
// (18, 21, 'sp4_v_b_22')
// (18, 22, 'sp4_v_b_11')

reg n57 = 0;
// (4, 17, 'neigh_op_tnr_5')
// (4, 18, 'neigh_op_rgt_5')
// (4, 18, 'sp12_h_r_1')
// (4, 19, 'neigh_op_bnr_5')
// (5, 17, 'neigh_op_top_5')
// (5, 18, 'local_g1_5')
// (5, 18, 'lutff_5/in_1')
// (5, 18, 'lutff_5/out')
// (5, 18, 'sp12_h_r_2')
// (5, 19, 'neigh_op_bot_5')
// (6, 17, 'neigh_op_tnl_5')
// (6, 18, 'neigh_op_lft_5')
// (6, 18, 'sp12_h_r_5')
// (6, 19, 'neigh_op_bnl_5')
// (7, 18, 'sp12_h_r_6')
// (8, 18, 'sp12_h_r_9')
// (9, 18, 'sp12_h_r_10')
// (10, 18, 'sp12_h_r_13')
// (10, 18, 'sp4_h_r_6')
// (11, 18, 'sp12_h_r_14')
// (11, 18, 'sp4_h_r_19')
// (12, 18, 'sp12_h_r_17')
// (12, 18, 'sp4_h_r_30')
// (13, 18, 'sp12_h_r_18')
// (13, 18, 'sp4_h_r_43')
// (14, 18, 'sp12_h_r_21')
// (14, 18, 'sp4_h_l_43')
// (14, 18, 'sp4_h_r_9')
// (15, 18, 'sp12_h_r_22')
// (15, 18, 'sp4_h_r_20')
// (16, 18, 'sp12_h_l_22')
// (16, 18, 'sp4_h_r_33')
// (17, 18, 'sp4_h_r_44')
// (17, 19, 'sp4_r_v_b_39')
// (17, 20, 'sp4_r_v_b_26')
// (17, 21, 'sp4_r_v_b_15')
// (17, 22, 'sp4_r_v_b_2')
// (18, 18, 'sp4_h_l_44')
// (18, 18, 'sp4_v_t_39')
// (18, 19, 'sp4_v_b_39')
// (18, 20, 'sp4_v_b_26')
// (18, 21, 'local_g1_7')
// (18, 21, 'lutff_4/in_0')
// (18, 21, 'sp4_v_b_15')
// (18, 22, 'sp4_v_b_2')

reg n58 = 0;
// (4, 17, 'neigh_op_tnr_6')
// (4, 18, 'neigh_op_rgt_6')
// (4, 19, 'neigh_op_bnr_6')
// (5, 12, 'sp12_v_t_23')
// (5, 13, 'sp12_v_b_23')
// (5, 14, 'sp12_v_b_20')
// (5, 15, 'sp12_v_b_19')
// (5, 16, 'sp12_v_b_16')
// (5, 17, 'neigh_op_top_6')
// (5, 17, 'sp12_v_b_15')
// (5, 18, 'local_g1_6')
// (5, 18, 'lutff_6/in_1')
// (5, 18, 'lutff_6/out')
// (5, 18, 'sp12_v_b_12')
// (5, 19, 'neigh_op_bot_6')
// (5, 19, 'sp12_v_b_11')
// (5, 20, 'sp12_v_b_8')
// (5, 21, 'sp12_v_b_7')
// (5, 22, 'sp12_v_b_4')
// (5, 23, 'sp12_v_b_3')
// (5, 24, 'sp12_h_r_0')
// (5, 24, 'sp12_v_b_0')
// (6, 17, 'neigh_op_tnl_6')
// (6, 18, 'neigh_op_lft_6')
// (6, 19, 'neigh_op_bnl_6')
// (6, 24, 'sp12_h_r_3')
// (7, 24, 'sp12_h_r_4')
// (8, 24, 'sp12_h_r_7')
// (9, 24, 'sp12_h_r_8')
// (10, 24, 'sp12_h_r_11')
// (11, 24, 'sp12_h_r_12')
// (12, 24, 'sp12_h_r_15')
// (13, 24, 'sp12_h_r_16')
// (14, 24, 'sp12_h_r_19')
// (14, 24, 'sp4_h_r_11')
// (15, 24, 'sp12_h_r_20')
// (15, 24, 'sp4_h_r_22')
// (16, 24, 'sp12_h_r_23')
// (16, 24, 'sp4_h_r_35')
// (17, 21, 'sp4_r_v_b_46')
// (17, 22, 'sp4_r_v_b_35')
// (17, 23, 'sp4_r_v_b_22')
// (17, 24, 'sp12_h_l_23')
// (17, 24, 'sp4_h_r_46')
// (17, 24, 'sp4_r_v_b_11')
// (18, 20, 'sp4_v_t_46')
// (18, 21, 'sp4_v_b_46')
// (18, 22, 'sp4_v_b_35')
// (18, 23, 'local_g0_6')
// (18, 23, 'lutff_6/in_0')
// (18, 23, 'sp4_v_b_22')
// (18, 24, 'sp4_h_l_46')
// (18, 24, 'sp4_v_b_11')

reg n59 = 0;
// (4, 17, 'sp12_h_r_1')
// (5, 17, 'sp12_h_r_2')
// (6, 17, 'sp12_h_r_5')
// (7, 17, 'sp12_h_r_6')
// (8, 17, 'sp12_h_r_9')
// (9, 17, 'local_g1_2')
// (9, 17, 'lutff_0/in_1')
// (9, 17, 'sp12_h_r_10')
// (10, 17, 'sp12_h_r_13')
// (11, 17, 'sp12_h_r_14')
// (11, 21, 'local_g0_2')
// (11, 21, 'lutff_3/in_1')
// (11, 21, 'sp4_h_r_10')
// (12, 17, 'sp12_h_r_17')
// (12, 21, 'sp4_h_r_23')
// (13, 17, 'sp12_h_r_18')
// (13, 21, 'sp4_h_r_34')
// (14, 17, 'sp12_h_r_21')
// (14, 18, 'sp4_r_v_b_40')
// (14, 19, 'sp4_r_v_b_29')
// (14, 20, 'sp4_r_v_b_16')
// (14, 21, 'sp4_h_r_47')
// (14, 21, 'sp4_r_v_b_5')
// (15, 11, 'neigh_op_tnr_5')
// (15, 12, 'neigh_op_rgt_5')
// (15, 12, 'sp12_h_r_1')
// (15, 12, 'sp12_v_t_22')
// (15, 12, 'sp4_r_v_b_42')
// (15, 13, 'neigh_op_bnr_5')
// (15, 13, 'sp12_v_b_22')
// (15, 13, 'sp4_r_v_b_31')
// (15, 14, 'sp12_v_b_21')
// (15, 14, 'sp4_r_v_b_18')
// (15, 15, 'sp12_v_b_18')
// (15, 15, 'sp4_r_v_b_7')
// (15, 16, 'local_g2_1')
// (15, 16, 'local_g3_1')
// (15, 16, 'lutff_1/in_1')
// (15, 16, 'lutff_2/in_2')
// (15, 16, 'lutff_3/in_3')
// (15, 16, 'lutff_4/in_3')
// (15, 16, 'lutff_5/in_0')
// (15, 16, 'lutff_6/in_1')
// (15, 16, 'lutff_7/in_1')
// (15, 16, 'sp12_v_b_17')
// (15, 17, 'sp12_h_r_22')
// (15, 17, 'sp12_v_b_14')
// (15, 17, 'sp4_v_t_40')
// (15, 18, 'sp12_v_b_13')
// (15, 18, 'sp4_v_b_40')
// (15, 19, 'sp12_v_b_10')
// (15, 19, 'sp4_v_b_29')
// (15, 20, 'sp12_v_b_9')
// (15, 20, 'sp4_v_b_16')
// (15, 21, 'sp12_v_b_6')
// (15, 21, 'sp4_h_l_47')
// (15, 21, 'sp4_v_b_5')
// (15, 22, 'sp12_v_b_5')
// (15, 23, 'sp12_v_b_2')
// (15, 24, 'sp12_v_b_1')
// (16, 5, 'sp12_v_t_22')
// (16, 6, 'sp12_v_b_22')
// (16, 7, 'sp12_v_b_21')
// (16, 8, 'sp12_v_b_18')
// (16, 9, 'sp12_v_b_17')
// (16, 10, 'sp12_v_b_14')
// (16, 11, 'neigh_op_top_5')
// (16, 11, 'sp12_v_b_13')
// (16, 11, 'sp4_v_t_42')
// (16, 12, 'local_g0_5')
// (16, 12, 'lutff_3/in_0')
// (16, 12, 'lutff_5/out')
// (16, 12, 'lutff_6/in_3')
// (16, 12, 'sp12_h_r_2')
// (16, 12, 'sp12_v_b_10')
// (16, 12, 'sp4_v_b_42')
// (16, 13, 'local_g0_5')
// (16, 13, 'lutff_2/in_3')
// (16, 13, 'lutff_4/in_3')
// (16, 13, 'lutff_6/in_3')
// (16, 13, 'neigh_op_bot_5')
// (16, 13, 'sp12_v_b_9')
// (16, 13, 'sp4_v_b_31')
// (16, 14, 'local_g0_2')
// (16, 14, 'local_g1_2')
// (16, 14, 'lutff_2/in_1')
// (16, 14, 'lutff_6/in_3')
// (16, 14, 'lutff_7/in_3')
// (16, 14, 'sp12_v_b_6')
// (16, 14, 'sp4_v_b_18')
// (16, 15, 'local_g0_7')
// (16, 15, 'lutff_1/in_0')
// (16, 15, 'lutff_2/in_3')
// (16, 15, 'lutff_4/in_3')
// (16, 15, 'lutff_5/in_0')
// (16, 15, 'lutff_7/in_0')
// (16, 15, 'sp12_v_b_5')
// (16, 15, 'sp4_v_b_7')
// (16, 16, 'sp12_v_b_2')
// (16, 17, 'sp12_h_l_22')
// (16, 17, 'sp12_v_b_1')
// (16, 17, 'sp12_v_t_22')
// (16, 18, 'sp12_v_b_22')
// (16, 19, 'sp12_v_b_21')
// (16, 20, 'local_g3_2')
// (16, 20, 'lutff_4/in_3')
// (16, 20, 'lutff_5/in_0')
// (16, 20, 'lutff_6/in_1')
// (16, 20, 'lutff_7/in_0')
// (16, 20, 'sp12_v_b_18')
// (16, 21, 'sp12_v_b_17')
// (16, 22, 'sp12_v_b_14')
// (16, 23, 'sp12_v_b_13')
// (16, 24, 'sp12_v_b_10')
// (16, 25, 'sp12_v_b_9')
// (16, 26, 'sp12_v_b_6')
// (16, 27, 'sp12_v_b_5')
// (16, 28, 'sp12_v_b_2')
// (16, 29, 'sp12_v_b_1')
// (17, 11, 'neigh_op_tnl_5')
// (17, 12, 'neigh_op_lft_5')
// (17, 12, 'sp12_h_r_5')
// (17, 13, 'neigh_op_bnl_5')
// (18, 12, 'sp12_h_r_6')
// (19, 12, 'local_g0_1')
// (19, 12, 'lutff_0/in_1')
// (19, 12, 'lutff_1/in_0')
// (19, 12, 'lutff_2/in_1')
// (19, 12, 'lutff_3/in_0')
// (19, 12, 'lutff_4/in_1')
// (19, 12, 'lutff_6/in_1')
// (19, 12, 'sp12_h_r_9')
// (20, 12, 'sp12_h_r_10')
// (21, 12, 'sp12_h_r_13')
// (22, 12, 'sp12_h_r_14')
// (22, 13, 'sp4_r_v_b_45')
// (22, 14, 'sp4_r_v_b_32')
// (22, 15, 'local_g3_5')
// (22, 15, 'lutff_0/in_0')
// (22, 15, 'lutff_1/in_3')
// (22, 15, 'lutff_2/in_0')
// (22, 15, 'lutff_3/in_3')
// (22, 15, 'lutff_4/in_0')
// (22, 15, 'lutff_5/in_3')
// (22, 15, 'lutff_6/in_0')
// (22, 15, 'lutff_7/in_3')
// (22, 15, 'sp4_r_v_b_21')
// (22, 16, 'sp4_r_v_b_8')
// (23, 12, 'sp12_h_r_17')
// (23, 12, 'sp4_h_r_8')
// (23, 12, 'sp4_v_t_45')
// (23, 13, 'sp4_v_b_45')
// (23, 14, 'sp4_v_b_32')
// (23, 15, 'sp4_v_b_21')
// (23, 16, 'sp4_v_b_8')
// (24, 12, 'sp12_h_r_18')
// (24, 12, 'sp4_h_r_21')
// (25, 12, 'sp12_h_r_21')
// (25, 12, 'sp4_h_r_32')
// (26, 12, 'sp12_h_r_22')
// (26, 12, 'sp4_h_r_45')
// (27, 12, 'sp12_h_l_22')
// (27, 12, 'sp4_h_l_45')

reg n60 = 0;
// (4, 18, 'neigh_op_tnr_0')
// (4, 18, 'sp4_r_v_b_45')
// (4, 19, 'neigh_op_rgt_0')
// (4, 19, 'sp4_r_v_b_32')
// (4, 20, 'neigh_op_bnr_0')
// (4, 20, 'sp4_r_v_b_21')
// (4, 21, 'sp4_r_v_b_8')
// (5, 17, 'sp4_v_t_45')
// (5, 18, 'neigh_op_top_0')
// (5, 18, 'sp4_v_b_45')
// (5, 19, 'local_g3_0')
// (5, 19, 'lutff_0/in_1')
// (5, 19, 'lutff_0/out')
// (5, 19, 'sp4_v_b_32')
// (5, 20, 'neigh_op_bot_0')
// (5, 20, 'sp4_v_b_21')
// (5, 21, 'sp4_h_r_2')
// (5, 21, 'sp4_v_b_8')
// (6, 18, 'neigh_op_tnl_0')
// (6, 19, 'neigh_op_lft_0')
// (6, 20, 'neigh_op_bnl_0')
// (6, 21, 'sp4_h_r_15')
// (7, 21, 'sp4_h_r_26')
// (8, 21, 'sp4_h_r_39')
// (9, 21, 'sp4_h_l_39')
// (9, 21, 'sp4_h_r_2')
// (10, 21, 'sp4_h_r_15')
// (11, 21, 'sp4_h_r_26')
// (12, 21, 'sp4_h_r_39')
// (13, 21, 'sp4_h_l_39')
// (13, 21, 'sp4_h_r_10')
// (14, 21, 'sp4_h_r_23')
// (15, 21, 'sp4_h_r_34')
// (16, 21, 'sp4_h_r_47')
// (17, 21, 'sp4_h_l_47')
// (17, 21, 'sp4_h_r_10')
// (18, 21, 'local_g0_7')
// (18, 21, 'lutff_0/in_1')
// (18, 21, 'sp4_h_r_23')
// (19, 21, 'sp4_h_r_34')
// (20, 21, 'sp4_h_r_47')
// (21, 21, 'sp4_h_l_47')

reg n61 = 0;
// (4, 18, 'neigh_op_tnr_1')
// (4, 18, 'sp4_r_v_b_47')
// (4, 19, 'neigh_op_rgt_1')
// (4, 19, 'sp4_r_v_b_34')
// (4, 20, 'neigh_op_bnr_1')
// (4, 20, 'sp4_r_v_b_23')
// (4, 21, 'sp4_r_v_b_10')
// (5, 17, 'sp4_v_t_47')
// (5, 18, 'neigh_op_top_1')
// (5, 18, 'sp4_v_b_47')
// (5, 19, 'local_g3_1')
// (5, 19, 'lutff_1/in_1')
// (5, 19, 'lutff_1/out')
// (5, 19, 'sp4_v_b_34')
// (5, 20, 'neigh_op_bot_1')
// (5, 20, 'sp4_v_b_23')
// (5, 21, 'sp4_h_r_4')
// (5, 21, 'sp4_v_b_10')
// (6, 18, 'neigh_op_tnl_1')
// (6, 19, 'neigh_op_lft_1')
// (6, 20, 'neigh_op_bnl_1')
// (6, 21, 'sp4_h_r_17')
// (7, 21, 'sp4_h_r_28')
// (8, 21, 'sp4_h_r_41')
// (9, 21, 'sp4_h_l_41')
// (9, 21, 'sp4_h_r_7')
// (10, 21, 'sp4_h_r_18')
// (11, 21, 'sp4_h_r_31')
// (12, 21, 'sp4_h_r_42')
// (13, 21, 'sp4_h_l_42')
// (13, 21, 'sp4_h_r_7')
// (14, 21, 'sp4_h_r_18')
// (15, 21, 'sp4_h_r_31')
// (16, 21, 'sp4_h_r_42')
// (17, 21, 'sp4_h_l_42')
// (17, 21, 'sp4_h_r_7')
// (18, 21, 'local_g0_2')
// (18, 21, 'lutff_1/in_3')
// (18, 21, 'sp4_h_r_18')
// (19, 21, 'sp4_h_r_31')
// (20, 21, 'sp4_h_r_42')
// (21, 21, 'sp4_h_l_42')

wire io_5_33_0;
// (4, 32, 'neigh_op_tnr_0')
// (4, 32, 'neigh_op_tnr_4')
// (5, 29, 'sp12_h_r_0')
// (5, 29, 'sp12_v_t_23')
// (5, 30, 'sp12_v_b_23')
// (5, 31, 'sp12_v_b_20')
// (5, 32, 'neigh_op_top_0')
// (5, 32, 'neigh_op_top_4')
// (5, 32, 'sp12_v_b_19')
// (5, 33, 'io_0/D_IN_0')
// (5, 33, 'io_0/PAD')
// (5, 33, 'span12_vert_16')
// (6, 29, 'sp12_h_r_3')
// (6, 32, 'neigh_op_tnl_0')
// (6, 32, 'neigh_op_tnl_4')
// (7, 29, 'sp12_h_r_4')
// (8, 29, 'sp12_h_r_7')
// (9, 29, 'sp12_h_r_8')
// (10, 29, 'sp12_h_r_11')
// (11, 29, 'sp12_h_r_12')
// (12, 29, 'sp12_h_r_15')
// (13, 29, 'sp12_h_r_16')
// (14, 29, 'sp12_h_r_19')
// (15, 29, 'sp12_h_r_20')
// (16, 22, 'sp4_r_v_b_41')
// (16, 23, 'sp4_r_v_b_28')
// (16, 24, 'local_g3_1')
// (16, 24, 'lutff_3/in_3')
// (16, 24, 'sp4_r_v_b_17')
// (16, 25, 'sp4_r_v_b_4')
// (16, 29, 'sp12_h_r_23')
// (17, 17, 'sp12_v_t_23')
// (17, 18, 'sp12_v_b_23')
// (17, 19, 'sp12_v_b_20')
// (17, 20, 'sp12_v_b_19')
// (17, 21, 'sp12_v_b_16')
// (17, 21, 'sp4_v_t_41')
// (17, 22, 'sp12_v_b_15')
// (17, 22, 'sp4_v_b_41')
// (17, 23, 'sp12_v_b_12')
// (17, 23, 'sp4_v_b_28')
// (17, 24, 'sp12_v_b_11')
// (17, 24, 'sp4_v_b_17')
// (17, 25, 'sp12_v_b_8')
// (17, 25, 'sp4_v_b_4')
// (17, 26, 'sp12_v_b_7')
// (17, 27, 'sp12_v_b_4')
// (17, 28, 'sp12_v_b_3')
// (17, 29, 'sp12_h_l_23')
// (17, 29, 'sp12_v_b_0')

wire io_6_0_1;
// (5, 0, 'span4_horz_r_3')
// (6, 0, 'io_1/D_OUT_0')
// (6, 0, 'io_1/PAD')
// (6, 0, 'local_g0_7')
// (6, 0, 'span4_horz_r_7')
// (7, 0, 'span4_horz_r_11')
// (8, 0, 'span4_horz_r_15')
// (8, 1, 'sp4_r_v_b_19')
// (8, 2, 'sp4_r_v_b_6')
// (8, 3, 'sp4_r_v_b_47')
// (8, 4, 'sp4_r_v_b_34')
// (8, 5, 'sp4_r_v_b_23')
// (8, 6, 'sp4_r_v_b_10')
// (8, 7, 'sp4_r_v_b_39')
// (8, 8, 'sp4_r_v_b_26')
// (8, 9, 'sp4_r_v_b_15')
// (8, 10, 'sp4_r_v_b_2')
// (9, 0, 'span4_horz_l_15')
// (9, 0, 'span4_vert_19')
// (9, 1, 'sp4_v_b_19')
// (9, 2, 'sp4_v_b_6')
// (9, 2, 'sp4_v_t_47')
// (9, 3, 'sp4_v_b_47')
// (9, 4, 'sp4_v_b_34')
// (9, 5, 'sp4_v_b_23')
// (9, 6, 'sp4_v_b_10')
// (9, 6, 'sp4_v_t_39')
// (9, 7, 'sp4_v_b_39')
// (9, 8, 'sp4_v_b_26')
// (9, 9, 'sp4_v_b_15')
// (9, 10, 'sp4_h_r_2')
// (9, 10, 'sp4_v_b_2')
// (10, 9, 'neigh_op_tnr_5')
// (10, 10, 'neigh_op_rgt_5')
// (10, 10, 'sp4_h_r_15')
// (10, 11, 'neigh_op_bnr_5')
// (11, 9, 'neigh_op_top_5')
// (11, 10, 'lutff_5/out')
// (11, 10, 'sp4_h_r_26')
// (11, 11, 'neigh_op_bot_5')
// (12, 9, 'neigh_op_tnl_5')
// (12, 10, 'neigh_op_lft_5')
// (12, 10, 'sp4_h_r_39')
// (12, 11, 'neigh_op_bnl_5')
// (13, 10, 'sp4_h_l_39')

wire n64;
// (5, 8, 'neigh_op_tnr_6')
// (5, 9, 'neigh_op_rgt_6')
// (5, 10, 'neigh_op_bnr_6')
// (6, 8, 'neigh_op_top_6')
// (6, 9, 'lutff_6/out')
// (6, 9, 'sp4_r_v_b_45')
// (6, 10, 'neigh_op_bot_6')
// (6, 10, 'sp4_r_v_b_32')
// (6, 11, 'sp4_r_v_b_21')
// (6, 12, 'local_g2_0')
// (6, 12, 'lutff_5/in_3')
// (6, 12, 'sp4_r_v_b_8')
// (7, 8, 'neigh_op_tnl_6')
// (7, 8, 'sp4_v_t_45')
// (7, 9, 'local_g1_6')
// (7, 9, 'lutff_6/in_3')
// (7, 9, 'neigh_op_lft_6')
// (7, 9, 'sp4_v_b_45')
// (7, 10, 'neigh_op_bnl_6')
// (7, 10, 'sp4_v_b_32')
// (7, 11, 'sp4_v_b_21')
// (7, 12, 'sp4_v_b_8')

reg n65 = 0;
// (5, 9, 'sp12_h_r_0')
// (6, 8, 'neigh_op_tnr_6')
// (6, 9, 'neigh_op_rgt_6')
// (6, 9, 'sp12_h_r_3')
// (6, 10, 'neigh_op_bnr_6')
// (7, 7, 'sp4_r_v_b_37')
// (7, 8, 'local_g0_6')
// (7, 8, 'lutff_5/in_3')
// (7, 8, 'neigh_op_top_6')
// (7, 8, 'sp4_r_v_b_24')
// (7, 9, 'local_g3_6')
// (7, 9, 'lutff_6/in_1')
// (7, 9, 'lutff_6/out')
// (7, 9, 'sp12_h_r_4')
// (7, 9, 'sp4_r_v_b_13')
// (7, 10, 'neigh_op_bot_6')
// (7, 10, 'sp4_r_v_b_0')
// (8, 6, 'sp4_v_t_37')
// (8, 7, 'sp4_v_b_37')
// (8, 8, 'neigh_op_tnl_6')
// (8, 8, 'sp4_v_b_24')
// (8, 9, 'neigh_op_lft_6')
// (8, 9, 'sp12_h_r_7')
// (8, 9, 'sp4_v_b_13')
// (8, 10, 'neigh_op_bnl_6')
// (8, 10, 'sp4_h_r_0')
// (8, 10, 'sp4_v_b_0')
// (9, 9, 'sp12_h_r_8')
// (9, 10, 'sp4_h_r_13')
// (10, 9, 'sp12_h_r_11')
// (10, 10, 'sp4_h_r_24')
// (11, 9, 'local_g1_4')
// (11, 9, 'lutff_4/in_3')
// (11, 9, 'lutff_5/in_0')
// (11, 9, 'sp12_h_r_12')
// (11, 10, 'local_g3_5')
// (11, 10, 'lutff_5/in_3')
// (11, 10, 'sp4_h_r_37')
// (12, 9, 'sp12_h_r_15')
// (12, 10, 'sp4_h_l_37')
// (13, 9, 'sp12_h_r_16')
// (14, 9, 'sp12_h_r_19')
// (15, 9, 'sp12_h_r_20')
// (16, 9, 'sp12_h_r_23')
// (17, 9, 'sp12_h_l_23')

wire n66;
// (5, 9, 'sp4_r_v_b_37')
// (5, 10, 'sp4_r_v_b_24')
// (5, 11, 'neigh_op_tnr_0')
// (5, 11, 'sp4_r_v_b_13')
// (5, 12, 'neigh_op_rgt_0')
// (5, 12, 'sp4_r_v_b_0')
// (5, 13, 'neigh_op_bnr_0')
// (6, 8, 'sp4_v_t_37')
// (6, 9, 'local_g2_5')
// (6, 9, 'lutff_6/in_3')
// (6, 9, 'sp4_v_b_37')
// (6, 10, 'sp4_v_b_24')
// (6, 11, 'neigh_op_top_0')
// (6, 11, 'sp4_v_b_13')
// (6, 12, 'lutff_0/out')
// (6, 12, 'sp4_h_r_0')
// (6, 12, 'sp4_v_b_0')
// (6, 13, 'neigh_op_bot_0')
// (7, 11, 'local_g3_0')
// (7, 11, 'lutff_1/in_0')
// (7, 11, 'lutff_6/in_3')
// (7, 11, 'neigh_op_tnl_0')
// (7, 12, 'local_g1_0')
// (7, 12, 'lutff_6/in_3')
// (7, 12, 'neigh_op_lft_0')
// (7, 12, 'sp4_h_r_13')
// (7, 13, 'neigh_op_bnl_0')
// (8, 12, 'sp4_h_r_24')
// (9, 12, 'local_g2_5')
// (9, 12, 'lutff_4/in_3')
// (9, 12, 'sp4_h_r_37')
// (10, 12, 'sp4_h_l_37')

reg n67 = 0;
// (5, 10, 'neigh_op_tnr_0')
// (5, 11, 'neigh_op_rgt_0')
// (5, 12, 'neigh_op_bnr_0')
// (6, 10, 'neigh_op_top_0')
// (6, 11, 'local_g3_0')
// (6, 11, 'lutff_0/in_1')
// (6, 11, 'lutff_0/out')
// (6, 12, 'local_g0_0')
// (6, 12, 'local_g1_0')
// (6, 12, 'lutff_0/in_0')
// (6, 12, 'lutff_2/in_1')
// (6, 12, 'neigh_op_bot_0')
// (7, 10, 'neigh_op_tnl_0')
// (7, 11, 'neigh_op_lft_0')
// (7, 12, 'neigh_op_bnl_0')

reg n68 = 0;
// (5, 10, 'neigh_op_tnr_1')
// (5, 11, 'neigh_op_rgt_1')
// (5, 12, 'neigh_op_bnr_1')
// (6, 10, 'neigh_op_top_1')
// (6, 11, 'local_g3_1')
// (6, 11, 'lutff_1/in_1')
// (6, 11, 'lutff_1/out')
// (6, 12, 'local_g1_1')
// (6, 12, 'lutff_1/in_3')
// (6, 12, 'lutff_2/in_0')
// (6, 12, 'neigh_op_bot_1')
// (7, 10, 'neigh_op_tnl_1')
// (7, 11, 'neigh_op_lft_1')
// (7, 12, 'neigh_op_bnl_1')

reg n69 = 0;
// (5, 10, 'neigh_op_tnr_2')
// (5, 11, 'neigh_op_rgt_2')
// (5, 12, 'neigh_op_bnr_2')
// (6, 10, 'neigh_op_top_2')
// (6, 11, 'local_g1_2')
// (6, 11, 'lutff_2/in_1')
// (6, 11, 'lutff_2/out')
// (6, 12, 'local_g0_2')
// (6, 12, 'lutff_0/in_2')
// (6, 12, 'lutff_2/in_2')
// (6, 12, 'neigh_op_bot_2')
// (7, 10, 'neigh_op_tnl_2')
// (7, 11, 'neigh_op_lft_2')
// (7, 12, 'neigh_op_bnl_2')

reg n70 = 0;
// (5, 10, 'neigh_op_tnr_3')
// (5, 11, 'neigh_op_rgt_3')
// (5, 12, 'neigh_op_bnr_3')
// (6, 10, 'neigh_op_top_3')
// (6, 11, 'local_g1_3')
// (6, 11, 'lutff_3/in_1')
// (6, 11, 'lutff_3/out')
// (6, 12, 'local_g0_3')
// (6, 12, 'local_g1_3')
// (6, 12, 'lutff_1/in_1')
// (6, 12, 'lutff_2/in_3')
// (6, 12, 'neigh_op_bot_3')
// (7, 10, 'neigh_op_tnl_3')
// (7, 11, 'neigh_op_lft_3')
// (7, 12, 'neigh_op_bnl_3')

reg n71 = 0;
// (5, 10, 'neigh_op_tnr_4')
// (5, 11, 'neigh_op_rgt_4')
// (5, 12, 'neigh_op_bnr_4')
// (6, 10, 'neigh_op_top_4')
// (6, 11, 'local_g3_4')
// (6, 11, 'lutff_4/in_1')
// (6, 11, 'lutff_4/out')
// (6, 12, 'local_g0_4')
// (6, 12, 'lutff_4/in_0')
// (6, 12, 'neigh_op_bot_4')
// (7, 10, 'neigh_op_tnl_4')
// (7, 11, 'neigh_op_lft_4')
// (7, 12, 'neigh_op_bnl_4')

reg n72 = 0;
// (5, 10, 'neigh_op_tnr_5')
// (5, 11, 'neigh_op_rgt_5')
// (5, 12, 'neigh_op_bnr_5')
// (6, 10, 'neigh_op_top_5')
// (6, 11, 'local_g1_5')
// (6, 11, 'lutff_5/in_1')
// (6, 11, 'lutff_5/out')
// (6, 12, 'local_g0_5')
// (6, 12, 'lutff_4/in_3')
// (6, 12, 'neigh_op_bot_5')
// (7, 10, 'neigh_op_tnl_5')
// (7, 11, 'neigh_op_lft_5')
// (7, 12, 'neigh_op_bnl_5')

reg n73 = 0;
// (5, 10, 'neigh_op_tnr_6')
// (5, 11, 'neigh_op_rgt_6')
// (5, 12, 'neigh_op_bnr_6')
// (6, 10, 'neigh_op_top_6')
// (6, 11, 'local_g1_6')
// (6, 11, 'lutff_6/in_1')
// (6, 11, 'lutff_6/out')
// (6, 12, 'local_g1_6')
// (6, 12, 'lutff_4/in_1')
// (6, 12, 'neigh_op_bot_6')
// (7, 10, 'neigh_op_tnl_6')
// (7, 11, 'neigh_op_lft_6')
// (7, 12, 'neigh_op_bnl_6')

reg n74 = 0;
// (5, 10, 'neigh_op_tnr_7')
// (5, 11, 'neigh_op_rgt_7')
// (5, 12, 'neigh_op_bnr_7')
// (6, 10, 'neigh_op_top_7')
// (6, 11, 'local_g2_7')
// (6, 11, 'lutff_7/in_0')
// (6, 11, 'lutff_7/out')
// (6, 12, 'local_g1_7')
// (6, 12, 'lutff_4/in_2')
// (6, 12, 'neigh_op_bot_7')
// (7, 10, 'neigh_op_tnl_7')
// (7, 11, 'neigh_op_lft_7')
// (7, 12, 'neigh_op_bnl_7')

reg n75 = 0;
// (5, 10, 'sp4_h_r_6')
// (5, 11, 'sp4_h_r_11')
// (6, 10, 'sp4_h_r_19')
// (6, 11, 'sp4_h_r_22')
// (6, 13, 'sp4_h_r_7')
// (7, 10, 'local_g2_6')
// (7, 10, 'lutff_7/in_3')
// (7, 10, 'sp4_h_r_30')
// (7, 11, 'local_g3_3')
// (7, 11, 'lutff_6/in_2')
// (7, 11, 'sp4_h_r_35')
// (7, 13, 'local_g1_2')
// (7, 13, 'lutff_5/in_2')
// (7, 13, 'sp4_h_r_18')
// (8, 10, 'sp4_h_r_43')
// (8, 11, 'neigh_op_tnr_7')
// (8, 11, 'sp4_h_r_46')
// (8, 11, 'sp4_r_v_b_43')
// (8, 12, 'neigh_op_rgt_7')
// (8, 12, 'sp4_r_v_b_30')
// (8, 12, 'sp4_r_v_b_46')
// (8, 13, 'neigh_op_bnr_7')
// (8, 13, 'sp4_h_r_31')
// (8, 13, 'sp4_r_v_b_19')
// (8, 13, 'sp4_r_v_b_35')
// (8, 14, 'sp4_r_v_b_22')
// (8, 14, 'sp4_r_v_b_6')
// (8, 15, 'sp4_r_v_b_11')
// (9, 10, 'local_g2_7')
// (9, 10, 'lutff_3/in_0')
// (9, 10, 'sp4_h_l_43')
// (9, 10, 'sp4_r_v_b_39')
// (9, 10, 'sp4_v_t_43')
// (9, 11, 'neigh_op_top_7')
// (9, 11, 'sp4_h_l_46')
// (9, 11, 'sp4_r_v_b_26')
// (9, 11, 'sp4_v_b_43')
// (9, 11, 'sp4_v_t_46')
// (9, 12, 'local_g1_7')
// (9, 12, 'lutff_2/in_2')
// (9, 12, 'lutff_7/in_1')
// (9, 12, 'lutff_7/out')
// (9, 12, 'sp4_r_v_b_15')
// (9, 12, 'sp4_v_b_30')
// (9, 12, 'sp4_v_b_46')
// (9, 13, 'neigh_op_bot_7')
// (9, 13, 'sp4_h_r_42')
// (9, 13, 'sp4_r_v_b_2')
// (9, 13, 'sp4_v_b_19')
// (9, 13, 'sp4_v_b_35')
// (9, 14, 'sp4_v_b_22')
// (9, 14, 'sp4_v_b_6')
// (9, 15, 'sp4_v_b_11')
// (10, 9, 'sp4_v_t_39')
// (10, 10, 'sp4_v_b_39')
// (10, 11, 'neigh_op_tnl_7')
// (10, 11, 'sp4_v_b_26')
// (10, 12, 'neigh_op_lft_7')
// (10, 12, 'sp4_v_b_15')
// (10, 13, 'neigh_op_bnl_7')
// (10, 13, 'sp4_h_l_42')
// (10, 13, 'sp4_v_b_2')

wire n76;
// (5, 11, 'neigh_op_tnr_1')
// (5, 12, 'neigh_op_rgt_1')
// (5, 13, 'neigh_op_bnr_1')
// (6, 11, 'neigh_op_top_1')
// (6, 12, 'local_g2_1')
// (6, 12, 'lutff_0/in_1')
// (6, 12, 'lutff_1/out')
// (6, 13, 'neigh_op_bot_1')
// (7, 11, 'neigh_op_tnl_1')
// (7, 12, 'neigh_op_lft_1')
// (7, 13, 'neigh_op_bnl_1')

wire n77;
// (5, 11, 'neigh_op_tnr_2')
// (5, 12, 'neigh_op_rgt_2')
// (5, 13, 'neigh_op_bnr_2')
// (6, 11, 'neigh_op_top_2')
// (6, 12, 'local_g2_2')
// (6, 12, 'lutff_2/out')
// (6, 12, 'lutff_5/in_1')
// (6, 13, 'neigh_op_bot_2')
// (7, 11, 'neigh_op_tnl_2')
// (7, 12, 'local_g1_2')
// (7, 12, 'lutff_2/in_1')
// (7, 12, 'neigh_op_lft_2')
// (7, 13, 'neigh_op_bnl_2')

wire n78;
// (5, 11, 'neigh_op_tnr_4')
// (5, 12, 'neigh_op_rgt_4')
// (5, 13, 'neigh_op_bnr_4')
// (6, 11, 'neigh_op_top_4')
// (6, 12, 'local_g1_4')
// (6, 12, 'lutff_0/in_3')
// (6, 12, 'lutff_4/out')
// (6, 13, 'neigh_op_bot_4')
// (7, 11, 'neigh_op_tnl_4')
// (7, 12, 'local_g1_4')
// (7, 12, 'lutff_2/in_3')
// (7, 12, 'neigh_op_lft_4')
// (7, 13, 'neigh_op_bnl_4')

reg n79 = 0;
// (5, 11, 'neigh_op_tnr_5')
// (5, 12, 'neigh_op_rgt_5')
// (5, 13, 'neigh_op_bnr_5')
// (6, 11, 'neigh_op_top_5')
// (6, 12, 'local_g2_5')
// (6, 12, 'lutff_5/in_0')
// (6, 12, 'lutff_5/out')
// (6, 13, 'neigh_op_bot_5')
// (7, 11, 'neigh_op_tnl_5')
// (7, 12, 'local_g1_5')
// (7, 12, 'lutff_2/in_0')
// (7, 12, 'neigh_op_lft_5')
// (7, 13, 'neigh_op_bnl_5')

wire n80;
// (5, 11, 'sp4_h_r_9')
// (5, 13, 'sp4_h_r_5')
// (6, 11, 'sp4_h_r_20')
// (6, 13, 'sp4_h_r_16')
// (7, 11, 'local_g2_1')
// (7, 11, 'lutff_6/in_1')
// (7, 11, 'sp4_h_r_33')
// (7, 13, 'local_g3_5')
// (7, 13, 'lutff_5/in_1')
// (7, 13, 'sp4_h_r_29')
// (8, 11, 'sp4_h_r_44')
// (8, 12, 'sp4_r_v_b_38')
// (8, 13, 'neigh_op_tnr_7')
// (8, 13, 'sp4_h_r_40')
// (8, 13, 'sp4_r_v_b_27')
// (8, 14, 'neigh_op_rgt_7')
// (8, 14, 'sp4_r_v_b_14')
// (8, 14, 'sp4_r_v_b_46')
// (8, 15, 'neigh_op_bnr_7')
// (8, 15, 'sp4_r_v_b_3')
// (8, 15, 'sp4_r_v_b_35')
// (8, 16, 'sp4_r_v_b_22')
// (8, 17, 'sp4_r_v_b_11')
// (9, 11, 'sp4_h_l_44')
// (9, 11, 'sp4_v_t_38')
// (9, 12, 'local_g3_6')
// (9, 12, 'lutff_2/in_3')
// (9, 12, 'lutff_7/in_0')
// (9, 12, 'sp4_v_b_38')
// (9, 13, 'neigh_op_top_7')
// (9, 13, 'sp4_h_l_40')
// (9, 13, 'sp4_v_b_27')
// (9, 13, 'sp4_v_t_46')
// (9, 14, 'lutff_7/out')
// (9, 14, 'sp4_v_b_14')
// (9, 14, 'sp4_v_b_46')
// (9, 15, 'neigh_op_bot_7')
// (9, 15, 'sp4_v_b_3')
// (9, 15, 'sp4_v_b_35')
// (9, 16, 'sp4_v_b_22')
// (9, 17, 'sp4_v_b_11')
// (10, 13, 'neigh_op_tnl_7')
// (10, 14, 'neigh_op_lft_7')
// (10, 15, 'neigh_op_bnl_7')

wire n81;
// (5, 11, 'sp4_r_v_b_46')
// (5, 12, 'neigh_op_tnr_3')
// (5, 12, 'sp4_r_v_b_35')
// (5, 13, 'neigh_op_rgt_3')
// (5, 13, 'sp4_r_v_b_22')
// (5, 14, 'neigh_op_bnr_3')
// (5, 14, 'sp4_r_v_b_11')
// (6, 10, 'sp4_v_t_46')
// (6, 11, 'local_g2_6')
// (6, 11, 'local_g3_6')
// (6, 11, 'lutff_0/in_0')
// (6, 11, 'lutff_1/in_0')
// (6, 11, 'lutff_2/in_0')
// (6, 11, 'lutff_3/in_0')
// (6, 11, 'lutff_4/in_0')
// (6, 11, 'lutff_5/in_0')
// (6, 11, 'lutff_6/in_0')
// (6, 11, 'lutff_7/in_1')
// (6, 11, 'sp4_v_b_46')
// (6, 12, 'neigh_op_top_3')
// (6, 12, 'sp4_v_b_35')
// (6, 13, 'lutff_3/out')
// (6, 13, 'sp4_v_b_22')
// (6, 14, 'neigh_op_bot_3')
// (6, 14, 'sp4_v_b_11')
// (7, 12, 'neigh_op_tnl_3')
// (7, 13, 'neigh_op_lft_3')
// (7, 14, 'neigh_op_bnl_3')

wire io_25_0_0;
// (5, 14, 'sp4_r_v_b_46')
// (5, 15, 'sp4_r_v_b_35')
// (5, 16, 'sp4_r_v_b_22')
// (5, 17, 'sp4_r_v_b_11')
// (6, 13, 'sp4_h_r_11')
// (6, 13, 'sp4_v_t_46')
// (6, 14, 'sp4_v_b_46')
// (6, 15, 'sp4_v_b_35')
// (6, 16, 'local_g0_6')
// (6, 16, 'lutff_0/in_0')
// (6, 16, 'sp4_v_b_22')
// (6, 17, 'sp4_v_b_11')
// (7, 13, 'sp4_h_r_22')
// (7, 14, 'sp4_r_v_b_47')
// (7, 15, 'sp4_r_v_b_34')
// (7, 16, 'local_g3_7')
// (7, 16, 'lutff_7/in_1')
// (7, 16, 'sp4_r_v_b_23')
// (7, 17, 'sp4_r_v_b_10')
// (8, 13, 'sp4_h_r_35')
// (8, 13, 'sp4_h_r_4')
// (8, 13, 'sp4_v_t_47')
// (8, 14, 'sp4_v_b_47')
// (8, 15, 'sp4_v_b_34')
// (8, 16, 'sp4_v_b_23')
// (8, 17, 'sp4_v_b_10')
// (9, 13, 'sp4_h_r_17')
// (9, 13, 'sp4_h_r_46')
// (9, 14, 'sp4_r_v_b_38')
// (9, 15, 'sp4_r_v_b_27')
// (9, 16, 'local_g2_6')
// (9, 16, 'lutff_3/in_3')
// (9, 16, 'lutff_4/in_0')
// (9, 16, 'sp4_r_v_b_14')
// (9, 17, 'sp4_r_v_b_3')
// (10, 13, 'sp4_h_l_46')
// (10, 13, 'sp4_h_r_28')
// (10, 13, 'sp4_h_r_3')
// (10, 13, 'sp4_v_t_38')
// (10, 14, 'sp4_v_b_38')
// (10, 15, 'sp4_v_b_27')
// (10, 16, 'sp4_v_b_14')
// (10, 17, 'sp4_v_b_3')
// (11, 13, 'sp4_h_r_14')
// (11, 13, 'sp4_h_r_41')
// (12, 13, 'sp4_h_l_41')
// (12, 13, 'sp4_h_r_1')
// (12, 13, 'sp4_h_r_27')
// (13, 13, 'sp12_h_r_0')
// (13, 13, 'sp4_h_r_12')
// (13, 13, 'sp4_h_r_38')
// (14, 13, 'sp12_h_r_3')
// (14, 13, 'sp4_h_l_38')
// (14, 13, 'sp4_h_r_25')
// (14, 13, 'sp4_h_r_3')
// (15, 13, 'sp12_h_r_4')
// (15, 13, 'sp4_h_r_14')
// (15, 13, 'sp4_h_r_36')
// (16, 13, 'sp12_h_r_7')
// (16, 13, 'sp4_h_l_36')
// (16, 13, 'sp4_h_r_27')
// (17, 13, 'sp12_h_r_8')
// (17, 13, 'sp4_h_r_38')
// (18, 13, 'sp12_h_r_11')
// (18, 13, 'sp4_h_l_38')
// (19, 13, 'sp12_h_r_12')
// (20, 13, 'sp12_h_r_15')
// (21, 13, 'sp12_h_r_16')
// (22, 13, 'sp12_h_r_19')
// (23, 13, 'sp12_h_r_20')
// (24, 1, 'neigh_op_bnr_0')
// (24, 1, 'neigh_op_bnr_4')
// (24, 13, 'sp12_h_r_23')
// (25, 0, 'io_0/D_IN_0')
// (25, 0, 'io_0/PAD')
// (25, 0, 'span12_vert_0')
// (25, 1, 'neigh_op_bot_0')
// (25, 1, 'neigh_op_bot_4')
// (25, 1, 'sp12_v_b_0')
// (25, 1, 'sp12_v_t_23')
// (25, 2, 'sp12_v_b_23')
// (25, 3, 'sp12_v_b_20')
// (25, 4, 'sp12_v_b_19')
// (25, 5, 'sp12_v_b_16')
// (25, 6, 'sp12_v_b_15')
// (25, 7, 'sp12_v_b_12')
// (25, 8, 'sp12_v_b_11')
// (25, 9, 'sp12_v_b_8')
// (25, 10, 'sp12_v_b_7')
// (25, 11, 'sp12_v_b_4')
// (25, 12, 'sp12_v_b_3')
// (25, 13, 'sp12_h_l_23')
// (25, 13, 'sp12_v_b_0')
// (26, 1, 'neigh_op_bnl_0')
// (26, 1, 'neigh_op_bnl_4')

wire n83;
// (5, 15, 'neigh_op_tnr_0')
// (5, 16, 'neigh_op_rgt_0')
// (5, 16, 'sp4_h_r_5')
// (5, 17, 'neigh_op_bnr_0')
// (6, 15, 'neigh_op_top_0')
// (6, 16, 'lutff_0/out')
// (6, 16, 'sp4_h_r_16')
// (6, 17, 'neigh_op_bot_0')
// (7, 15, 'neigh_op_tnl_0')
// (7, 16, 'neigh_op_lft_0')
// (7, 16, 'sp4_h_r_29')
// (7, 17, 'neigh_op_bnl_0')
// (8, 16, 'sp4_h_r_40')
// (9, 16, 'sp4_h_l_40')
// (9, 16, 'sp4_h_r_8')
// (10, 16, 'sp4_h_r_21')
// (11, 16, 'local_g2_0')
// (11, 16, 'lutff_4/in_2')
// (11, 16, 'sp4_h_r_32')
// (12, 16, 'sp4_h_r_45')
// (13, 16, 'sp4_h_l_45')

reg n84 = 0;
// (5, 15, 'sp4_h_r_2')
// (6, 15, 'sp4_h_r_15')
// (7, 15, 'local_g3_2')
// (7, 15, 'lutff_2/in_1')
// (7, 15, 'sp4_h_r_26')
// (8, 12, 'sp4_r_v_b_44')
// (8, 13, 'neigh_op_tnr_2')
// (8, 13, 'sp4_r_v_b_33')
// (8, 14, 'neigh_op_rgt_2')
// (8, 14, 'sp4_r_v_b_20')
// (8, 15, 'neigh_op_bnr_2')
// (8, 15, 'sp4_h_r_39')
// (8, 15, 'sp4_r_v_b_9')
// (9, 11, 'sp4_v_t_44')
// (9, 12, 'sp4_v_b_44')
// (9, 13, 'neigh_op_top_2')
// (9, 13, 'sp4_v_b_33')
// (9, 14, 'local_g2_2')
// (9, 14, 'lutff_2/in_2')
// (9, 14, 'lutff_2/out')
// (9, 14, 'sp4_v_b_20')
// (9, 15, 'neigh_op_bot_2')
// (9, 15, 'sp4_h_l_39')
// (9, 15, 'sp4_v_b_9')
// (10, 13, 'neigh_op_tnl_2')
// (10, 14, 'neigh_op_lft_2')
// (10, 15, 'neigh_op_bnl_2')

wire n85;
// (5, 17, 'carry_in_mux')
// (5, 17, 'lutff_0/in_3')

wire n86;
// (5, 17, 'lutff_0/cout')
// (5, 17, 'lutff_1/in_3')

wire n87;
// (5, 17, 'lutff_1/cout')
// (5, 17, 'lutff_2/in_3')

wire n88;
// (5, 17, 'lutff_2/cout')
// (5, 17, 'lutff_3/in_3')

wire n89;
// (5, 17, 'lutff_3/cout')
// (5, 17, 'lutff_4/in_3')

wire n90;
// (5, 17, 'lutff_4/cout')
// (5, 17, 'lutff_5/in_3')

wire n91;
// (5, 17, 'lutff_5/cout')
// (5, 17, 'lutff_6/in_3')

wire n92;
// (5, 17, 'lutff_6/cout')
// (5, 17, 'lutff_7/in_3')

wire n93;
// (5, 17, 'lutff_7/cout')
// (5, 18, 'carry_in')
// (5, 18, 'carry_in_mux')
// (5, 18, 'lutff_0/in_3')

wire n94;
// (5, 18, 'lutff_0/cout')
// (5, 18, 'lutff_1/in_3')

wire n95;
// (5, 18, 'lutff_1/cout')
// (5, 18, 'lutff_2/in_3')

wire n96;
// (5, 18, 'lutff_2/cout')
// (5, 18, 'lutff_3/in_3')

wire n97;
// (5, 18, 'lutff_3/cout')
// (5, 18, 'lutff_4/in_3')

wire n98;
// (5, 18, 'lutff_4/cout')
// (5, 18, 'lutff_5/in_3')

wire n99;
// (5, 18, 'lutff_5/cout')
// (5, 18, 'lutff_6/in_3')

wire n100;
// (5, 18, 'lutff_6/cout')
// (5, 18, 'lutff_7/in_3')

wire n101;
// (5, 18, 'lutff_7/cout')
// (5, 19, 'carry_in')
// (5, 19, 'carry_in_mux')
// (5, 19, 'lutff_0/in_3')

wire n102;
// (5, 19, 'lutff_0/cout')
// (5, 19, 'lutff_1/in_3')

wire n103;
// (5, 19, 'lutff_1/cout')
// (5, 19, 'lutff_2/in_3')

reg n104 = 0;
// (5, 23, 'sp12_h_r_1')
// (6, 23, 'sp12_h_r_2')
// (7, 23, 'sp12_h_r_5')
// (8, 23, 'sp12_h_r_6')
// (9, 23, 'sp12_h_r_9')
// (10, 23, 'sp12_h_r_10')
// (11, 23, 'sp12_h_r_13')
// (12, 23, 'sp12_h_r_14')
// (13, 23, 'sp12_h_r_17')
// (14, 23, 'sp12_h_r_18')
// (15, 22, 'neigh_op_tnr_7')
// (15, 23, 'neigh_op_rgt_7')
// (15, 23, 'sp12_h_r_21')
// (15, 24, 'neigh_op_bnr_7')
// (16, 22, 'neigh_op_top_7')
// (16, 23, 'lutff_7/out')
// (16, 23, 'sp12_h_r_22')
// (16, 24, 'neigh_op_bot_7')
// (17, 22, 'neigh_op_tnl_7')
// (17, 23, 'neigh_op_lft_7')
// (17, 23, 'sp12_h_l_22')
// (17, 23, 'sp12_h_r_1')
// (17, 24, 'neigh_op_bnl_7')
// (18, 23, 'sp12_h_r_2')
// (19, 23, 'sp12_h_r_5')
// (20, 23, 'sp12_h_r_6')
// (21, 23, 'sp12_h_r_9')
// (22, 23, 'sp12_h_r_10')
// (23, 23, 'sp12_h_r_13')
// (24, 23, 'sp12_h_r_14')
// (25, 23, 'sp12_h_r_17')
// (26, 23, 'sp12_h_r_18')
// (27, 23, 'sp12_h_r_21')
// (28, 23, 'sp12_h_r_22')
// (29, 23, 'sp12_h_l_22')
// (29, 23, 'sp12_v_t_22')
// (29, 24, 'sp12_v_b_22')
// (29, 25, 'sp12_v_b_21')
// (29, 26, 'sp12_v_b_18')
// (29, 27, 'sp12_v_b_17')
// (29, 28, 'sp12_v_b_14')
// (29, 29, 'sp12_v_b_13')
// (29, 30, 'sp12_v_b_10')
// (29, 31, 'sp12_v_b_9')
// (29, 32, 'sp12_v_b_6')
// (29, 33, 'io_0/D_OUT_0')
// (29, 33, 'local_g1_5')
// (29, 33, 'span12_vert_5')

wire io_6_33_0;
// (5, 32, 'neigh_op_tnr_0')
// (5, 32, 'neigh_op_tnr_4')
// (6, 25, 'sp12_h_r_0')
// (6, 25, 'sp12_v_t_23')
// (6, 26, 'sp12_v_b_23')
// (6, 27, 'sp12_v_b_20')
// (6, 28, 'sp12_v_b_19')
// (6, 29, 'sp12_v_b_16')
// (6, 30, 'sp12_v_b_15')
// (6, 31, 'sp12_v_b_12')
// (6, 32, 'neigh_op_top_0')
// (6, 32, 'neigh_op_top_4')
// (6, 32, 'sp12_v_b_11')
// (6, 33, 'io_0/D_IN_0')
// (6, 33, 'io_0/PAD')
// (6, 33, 'span12_vert_8')
// (7, 25, 'sp12_h_r_3')
// (7, 32, 'neigh_op_tnl_0')
// (7, 32, 'neigh_op_tnl_4')
// (8, 25, 'sp12_h_r_4')
// (9, 25, 'sp12_h_r_7')
// (10, 25, 'sp12_h_r_8')
// (11, 25, 'sp12_h_r_11')
// (12, 25, 'sp12_h_r_12')
// (13, 25, 'sp12_h_r_15')
// (13, 25, 'sp4_h_r_9')
// (14, 25, 'sp12_h_r_16')
// (14, 25, 'sp4_h_r_20')
// (15, 25, 'sp12_h_r_19')
// (15, 25, 'sp4_h_r_33')
// (16, 22, 'sp4_r_v_b_38')
// (16, 23, 'sp4_r_v_b_27')
// (16, 24, 'local_g2_6')
// (16, 24, 'lutff_2/in_0')
// (16, 24, 'sp4_r_v_b_14')
// (16, 25, 'sp12_h_r_20')
// (16, 25, 'sp4_h_r_44')
// (16, 25, 'sp4_r_v_b_3')
// (17, 21, 'sp4_v_t_38')
// (17, 22, 'sp4_v_b_38')
// (17, 23, 'sp4_v_b_27')
// (17, 24, 'sp4_v_b_14')
// (17, 25, 'sp12_h_r_23')
// (17, 25, 'sp4_h_l_44')
// (17, 25, 'sp4_v_b_3')
// (18, 25, 'sp12_h_l_23')

wire io_6_33_1;
// (5, 32, 'neigh_op_tnr_2')
// (5, 32, 'neigh_op_tnr_6')
// (6, 27, 'sp12_h_r_0')
// (6, 27, 'sp12_v_t_23')
// (6, 28, 'sp12_v_b_23')
// (6, 29, 'sp12_v_b_20')
// (6, 30, 'sp12_v_b_19')
// (6, 31, 'sp12_v_b_16')
// (6, 32, 'neigh_op_top_2')
// (6, 32, 'neigh_op_top_6')
// (6, 32, 'sp12_v_b_15')
// (6, 33, 'io_1/D_IN_0')
// (6, 33, 'io_1/PAD')
// (6, 33, 'span12_vert_12')
// (7, 27, 'sp12_h_r_3')
// (7, 32, 'neigh_op_tnl_2')
// (7, 32, 'neigh_op_tnl_6')
// (8, 27, 'sp12_h_r_4')
// (9, 27, 'sp12_h_r_7')
// (10, 27, 'sp12_h_r_8')
// (11, 27, 'sp12_h_r_11')
// (12, 27, 'sp12_h_r_12')
// (13, 27, 'sp12_h_r_15')
// (13, 27, 'sp4_h_r_9')
// (14, 27, 'sp12_h_r_16')
// (14, 27, 'sp4_h_r_20')
// (15, 27, 'sp12_h_r_19')
// (15, 27, 'sp4_h_r_33')
// (16, 24, 'local_g3_4')
// (16, 24, 'lutff_1/in_0')
// (16, 24, 'sp4_r_v_b_44')
// (16, 25, 'sp4_r_v_b_33')
// (16, 26, 'sp4_r_v_b_20')
// (16, 27, 'sp12_h_r_20')
// (16, 27, 'sp4_h_r_44')
// (16, 27, 'sp4_r_v_b_9')
// (17, 23, 'sp4_v_t_44')
// (17, 24, 'sp4_v_b_44')
// (17, 25, 'sp4_v_b_33')
// (17, 26, 'sp4_v_b_20')
// (17, 27, 'sp12_h_r_23')
// (17, 27, 'sp4_h_l_44')
// (17, 27, 'sp4_v_b_9')
// (18, 27, 'sp12_h_l_23')

reg n107 = 0;
// (6, 9, 'local_g2_4')
// (6, 9, 'lutff_6/in_0')
// (6, 9, 'sp4_r_v_b_36')
// (6, 10, 'neigh_op_tnr_6')
// (6, 10, 'sp4_r_v_b_25')
// (6, 11, 'neigh_op_rgt_6')
// (6, 11, 'sp4_r_v_b_12')
// (6, 12, 'neigh_op_bnr_6')
// (6, 12, 'sp4_r_v_b_1')
// (7, 8, 'sp4_v_t_36')
// (7, 9, 'sp4_v_b_36')
// (7, 10, 'neigh_op_top_6')
// (7, 10, 'sp4_v_b_25')
// (7, 11, 'local_g2_6')
// (7, 11, 'lutff_6/in_0')
// (7, 11, 'lutff_6/out')
// (7, 11, 'sp4_v_b_12')
// (7, 12, 'local_g1_6')
// (7, 12, 'lutff_6/in_1')
// (7, 12, 'neigh_op_bot_6')
// (7, 12, 'sp4_v_b_1')
// (8, 10, 'neigh_op_tnl_6')
// (8, 11, 'neigh_op_lft_6')
// (8, 12, 'neigh_op_bnl_6')

reg n108 = 0;
// (6, 9, 'neigh_op_tnr_3')
// (6, 10, 'neigh_op_rgt_3')
// (6, 10, 'sp4_h_r_11')
// (6, 11, 'neigh_op_bnr_3')
// (7, 9, 'local_g1_3')
// (7, 9, 'lutff_6/in_2')
// (7, 9, 'neigh_op_top_3')
// (7, 10, 'local_g0_3')
// (7, 10, 'lutff_3/in_0')
// (7, 10, 'lutff_3/out')
// (7, 10, 'sp4_h_r_22')
// (7, 10, 'sp4_r_v_b_39')
// (7, 11, 'local_g0_3')
// (7, 11, 'lutff_1/in_2')
// (7, 11, 'neigh_op_bot_3')
// (7, 11, 'sp4_r_v_b_26')
// (7, 12, 'local_g2_7')
// (7, 12, 'lutff_7/in_0')
// (7, 12, 'sp4_r_v_b_15')
// (7, 13, 'sp4_r_v_b_2')
// (8, 9, 'neigh_op_tnl_3')
// (8, 9, 'sp4_v_t_39')
// (8, 10, 'neigh_op_lft_3')
// (8, 10, 'sp4_h_r_35')
// (8, 10, 'sp4_v_b_39')
// (8, 11, 'neigh_op_bnl_3')
// (8, 11, 'sp4_v_b_26')
// (8, 12, 'sp4_v_b_15')
// (8, 13, 'sp4_v_b_2')
// (9, 10, 'sp4_h_r_46')
// (9, 11, 'sp4_r_v_b_46')
// (9, 12, 'local_g2_3')
// (9, 12, 'lutff_1/in_2')
// (9, 12, 'lutff_2/in_1')
// (9, 12, 'sp4_r_v_b_35')
// (9, 13, 'sp4_r_v_b_22')
// (9, 14, 'sp4_r_v_b_11')
// (10, 10, 'sp4_h_l_46')
// (10, 10, 'sp4_v_t_46')
// (10, 11, 'sp4_v_b_46')
// (10, 12, 'sp4_v_b_35')
// (10, 13, 'sp4_v_b_22')
// (10, 14, 'sp4_v_b_11')

reg n109 = 0;
// (6, 9, 'neigh_op_tnr_6')
// (6, 10, 'neigh_op_rgt_6')
// (6, 11, 'neigh_op_bnr_6')
// (7, 9, 'local_g0_6')
// (7, 9, 'lutff_6/in_0')
// (7, 9, 'neigh_op_top_6')
// (7, 9, 'sp4_r_v_b_40')
// (7, 10, 'local_g0_6')
// (7, 10, 'lutff_3/in_1')
// (7, 10, 'lutff_6/out')
// (7, 10, 'sp4_r_v_b_29')
// (7, 10, 'sp4_r_v_b_45')
// (7, 11, 'local_g0_6')
// (7, 11, 'lutff_1/in_1')
// (7, 11, 'neigh_op_bot_6')
// (7, 11, 'sp4_r_v_b_16')
// (7, 11, 'sp4_r_v_b_32')
// (7, 12, 'local_g3_5')
// (7, 12, 'lutff_7/in_1')
// (7, 12, 'sp4_r_v_b_21')
// (7, 12, 'sp4_r_v_b_5')
// (7, 13, 'sp4_r_v_b_8')
// (8, 8, 'sp4_v_t_40')
// (8, 9, 'neigh_op_tnl_6')
// (8, 9, 'sp4_v_b_40')
// (8, 9, 'sp4_v_t_45')
// (8, 10, 'neigh_op_lft_6')
// (8, 10, 'sp4_v_b_29')
// (8, 10, 'sp4_v_b_45')
// (8, 11, 'neigh_op_bnl_6')
// (8, 11, 'sp4_v_b_16')
// (8, 11, 'sp4_v_b_32')
// (8, 12, 'sp4_h_r_5')
// (8, 12, 'sp4_v_b_21')
// (8, 12, 'sp4_v_b_5')
// (8, 13, 'sp4_v_b_8')
// (9, 12, 'local_g0_0')
// (9, 12, 'lutff_2/in_0')
// (9, 12, 'sp4_h_r_16')
// (10, 12, 'sp4_h_r_29')
// (11, 12, 'sp4_h_r_40')
// (12, 12, 'sp4_h_l_40')

reg n110 = 0;
// (6, 9, 'sp4_r_v_b_42')
// (6, 10, 'neigh_op_tnr_1')
// (6, 10, 'sp4_r_v_b_31')
// (6, 11, 'neigh_op_rgt_1')
// (6, 11, 'sp4_r_v_b_18')
// (6, 12, 'neigh_op_bnr_1')
// (6, 12, 'sp4_r_v_b_7')
// (7, 8, 'sp4_v_t_42')
// (7, 9, 'sp4_v_b_42')
// (7, 10, 'neigh_op_top_1')
// (7, 10, 'sp4_v_b_31')
// (7, 11, 'local_g3_1')
// (7, 11, 'lutff_1/in_3')
// (7, 11, 'lutff_1/out')
// (7, 11, 'sp4_v_b_18')
// (7, 12, 'local_g1_1')
// (7, 12, 'lutff_6/in_0')
// (7, 12, 'neigh_op_bot_1')
// (7, 12, 'sp4_h_r_1')
// (7, 12, 'sp4_v_b_7')
// (8, 10, 'neigh_op_tnl_1')
// (8, 11, 'neigh_op_lft_1')
// (8, 12, 'neigh_op_bnl_1')
// (8, 12, 'sp4_h_r_12')
// (9, 12, 'local_g2_1')
// (9, 12, 'lutff_4/in_1')
// (9, 12, 'sp4_h_r_25')
// (10, 12, 'sp4_h_r_36')
// (11, 12, 'sp4_h_l_36')

wire n111;
// (6, 10, 'sp4_r_v_b_44')
// (6, 11, 'neigh_op_tnr_2')
// (6, 11, 'sp4_r_v_b_33')
// (6, 12, 'neigh_op_rgt_2')
// (6, 12, 'sp4_r_v_b_20')
// (6, 13, 'neigh_op_bnr_2')
// (6, 13, 'sp4_r_v_b_9')
// (7, 9, 'sp4_v_t_44')
// (7, 10, 'local_g2_4')
// (7, 10, 'lutff_3/in_3')
// (7, 10, 'sp4_v_b_44')
// (7, 11, 'neigh_op_top_2')
// (7, 11, 'sp4_v_b_33')
// (7, 12, 'local_g2_2')
// (7, 12, 'lutff_2/out')
// (7, 12, 'lutff_7/in_3')
// (7, 12, 'sp4_v_b_20')
// (7, 13, 'neigh_op_bot_2')
// (7, 13, 'sp4_v_b_9')
// (8, 11, 'neigh_op_tnl_2')
// (8, 12, 'neigh_op_lft_2')
// (8, 13, 'neigh_op_bnl_2')

wire n112;
// (6, 11, 'carry_in_mux')
// (6, 11, 'lutff_0/in_3')

wire n113;
// (6, 11, 'lutff_0/cout')
// (6, 11, 'lutff_1/in_3')

wire n114;
// (6, 11, 'lutff_1/cout')
// (6, 11, 'lutff_2/in_3')

wire n115;
// (6, 11, 'lutff_2/cout')
// (6, 11, 'lutff_3/in_3')

wire n116;
// (6, 11, 'lutff_3/cout')
// (6, 11, 'lutff_4/in_3')

wire n117;
// (6, 11, 'lutff_4/cout')
// (6, 11, 'lutff_5/in_3')

wire n118;
// (6, 11, 'lutff_5/cout')
// (6, 11, 'lutff_6/in_3')

wire n119;
// (6, 11, 'lutff_6/cout')
// (6, 11, 'lutff_7/in_3')

wire n120;
// (6, 11, 'neigh_op_tnr_5')
// (6, 12, 'neigh_op_rgt_5')
// (6, 12, 'sp4_r_v_b_42')
// (6, 13, 'neigh_op_bnr_5')
// (6, 13, 'sp4_r_v_b_31')
// (6, 14, 'sp4_r_v_b_18')
// (6, 15, 'sp4_r_v_b_7')
// (7, 11, 'neigh_op_top_5')
// (7, 11, 'sp4_h_r_7')
// (7, 11, 'sp4_v_t_42')
// (7, 12, 'lutff_5/out')
// (7, 12, 'sp4_h_r_10')
// (7, 12, 'sp4_v_b_42')
// (7, 13, 'neigh_op_bot_5')
// (7, 13, 'sp4_v_b_31')
// (7, 14, 'sp4_v_b_18')
// (7, 15, 'sp4_v_b_7')
// (8, 11, 'neigh_op_tnl_5')
// (8, 11, 'sp4_h_r_18')
// (8, 12, 'neigh_op_lft_5')
// (8, 12, 'sp4_h_r_23')
// (8, 13, 'neigh_op_bnl_5')
// (9, 11, 'sp4_h_r_31')
// (9, 12, 'sp4_h_r_34')
// (10, 11, 'sp4_h_r_42')
// (10, 12, 'sp4_h_r_47')
// (10, 12, 'sp4_r_v_b_42')
// (10, 13, 'local_g0_7')
// (10, 13, 'local_g3_7')
// (10, 13, 'lutff_0/in_0')
// (10, 13, 'lutff_1/in_0')
// (10, 13, 'lutff_2/in_0')
// (10, 13, 'lutff_3/in_0')
// (10, 13, 'lutff_4/in_0')
// (10, 13, 'lutff_5/in_0')
// (10, 13, 'lutff_6/in_0')
// (10, 13, 'lutff_7/in_1')
// (10, 13, 'sp4_r_v_b_31')
// (10, 13, 'sp4_r_v_b_47')
// (10, 14, 'sp4_r_v_b_18')
// (10, 14, 'sp4_r_v_b_34')
// (10, 15, 'sp4_r_v_b_23')
// (10, 15, 'sp4_r_v_b_7')
// (10, 16, 'sp4_r_v_b_10')
// (11, 11, 'sp4_h_l_42')
// (11, 11, 'sp4_v_t_42')
// (11, 12, 'sp4_h_l_47')
// (11, 12, 'sp4_v_b_42')
// (11, 12, 'sp4_v_t_47')
// (11, 13, 'sp4_v_b_31')
// (11, 13, 'sp4_v_b_47')
// (11, 14, 'sp4_v_b_18')
// (11, 14, 'sp4_v_b_34')
// (11, 15, 'sp4_v_b_23')
// (11, 15, 'sp4_v_b_7')
// (11, 16, 'sp4_v_b_10')

wire n121;
// (6, 11, 'neigh_op_tnr_6')
// (6, 12, 'neigh_op_rgt_6')
// (6, 12, 'sp4_h_r_1')
// (6, 13, 'neigh_op_bnr_6')
// (7, 11, 'neigh_op_top_6')
// (7, 12, 'lutff_6/out')
// (7, 12, 'sp4_h_r_12')
// (7, 13, 'neigh_op_bot_6')
// (8, 11, 'neigh_op_tnl_6')
// (8, 12, 'neigh_op_lft_6')
// (8, 12, 'sp4_h_r_25')
// (8, 13, 'neigh_op_bnl_6')
// (9, 12, 'local_g2_4')
// (9, 12, 'lutff_1/in_1')
// (9, 12, 'sp4_h_r_36')
// (10, 12, 'sp4_h_l_36')

wire n122;
// (6, 11, 'neigh_op_tnr_7')
// (6, 12, 'neigh_op_rgt_7')
// (6, 13, 'neigh_op_bnr_7')
// (7, 11, 'neigh_op_top_7')
// (7, 12, 'lutff_7/out')
// (7, 13, 'local_g1_7')
// (7, 13, 'lutff_5/in_3')
// (7, 13, 'neigh_op_bot_7')
// (8, 11, 'neigh_op_tnl_7')
// (8, 12, 'neigh_op_lft_7')
// (8, 13, 'neigh_op_bnl_7')

wire n123;
// (6, 12, 'lutff_4/lout')
// (6, 12, 'lutff_5/in_2')

reg n124 = 0;
// (6, 12, 'neigh_op_tnr_5')
// (6, 13, 'local_g3_5')
// (6, 13, 'lutff_3/in_3')
// (6, 13, 'neigh_op_rgt_5')
// (6, 14, 'neigh_op_bnr_5')
// (7, 12, 'neigh_op_top_5')
// (7, 13, 'local_g2_5')
// (7, 13, 'lutff_5/in_0')
// (7, 13, 'lutff_5/out')
// (7, 14, 'neigh_op_bot_5')
// (8, 12, 'neigh_op_tnl_5')
// (8, 13, 'neigh_op_lft_5')
// (8, 14, 'neigh_op_bnl_5')

reg n125 = 0;
// (6, 12, 'sp12_h_r_1')
// (7, 12, 'local_g0_2')
// (7, 12, 'lutff_1/in_1')
// (7, 12, 'sp12_h_r_2')
// (8, 12, 'sp12_h_r_5')
// (9, 12, 'sp12_h_r_6')
// (10, 12, 'sp12_h_r_9')
// (11, 12, 'sp12_h_r_10')
// (12, 12, 'sp12_h_r_13')
// (13, 12, 'sp12_h_r_14')
// (14, 11, 'neigh_op_tnr_5')
// (14, 12, 'neigh_op_rgt_5')
// (14, 12, 'sp12_h_r_17')
// (14, 13, 'neigh_op_bnr_5')
// (15, 11, 'neigh_op_top_5')
// (15, 12, 'local_g1_5')
// (15, 12, 'lutff_5/out')
// (15, 12, 'lutff_7/in_3')
// (15, 12, 'sp12_h_r_18')
// (15, 13, 'neigh_op_bot_5')
// (16, 11, 'neigh_op_tnl_5')
// (16, 12, 'neigh_op_lft_5')
// (16, 12, 'sp12_h_r_21')
// (16, 13, 'neigh_op_bnl_5')
// (17, 12, 'sp12_h_r_22')
// (18, 12, 'sp12_h_l_22')

reg n126 = 0;
// (6, 13, 'sp4_r_v_b_37')
// (6, 14, 'sp4_r_v_b_24')
// (6, 15, 'sp4_r_v_b_13')
// (6, 16, 'sp4_r_v_b_0')
// (7, 12, 'sp4_h_r_0')
// (7, 12, 'sp4_v_t_37')
// (7, 13, 'sp4_v_b_37')
// (7, 14, 'sp4_v_b_24')
// (7, 15, 'local_g0_5')
// (7, 15, 'lutff_2/in_3')
// (7, 15, 'sp4_v_b_13')
// (7, 16, 'sp4_v_b_0')
// (8, 12, 'sp4_h_r_13')
// (9, 12, 'sp4_h_r_24')
// (10, 12, 'sp4_h_r_37')
// (11, 12, 'sp4_h_l_37')
// (11, 12, 'sp4_h_r_0')
// (12, 12, 'sp4_h_r_13')
// (13, 12, 'sp4_h_r_24')
// (14, 11, 'neigh_op_tnr_0')
// (14, 12, 'neigh_op_rgt_0')
// (14, 12, 'sp4_h_r_37')
// (14, 13, 'neigh_op_bnr_0')
// (15, 11, 'neigh_op_top_0')
// (15, 12, 'local_g0_0')
// (15, 12, 'lutff_0/in_2')
// (15, 12, 'lutff_0/out')
// (15, 12, 'sp4_h_l_37')
// (15, 12, 'sp4_h_r_0')
// (15, 13, 'neigh_op_bot_0')
// (16, 11, 'neigh_op_tnl_0')
// (16, 12, 'neigh_op_lft_0')
// (16, 12, 'sp4_h_r_13')
// (16, 13, 'neigh_op_bnl_0')
// (17, 12, 'sp4_h_r_24')
// (18, 12, 'sp4_h_r_37')
// (19, 12, 'sp4_h_l_37')

wire n127;
// (6, 14, 'sp12_h_r_0')
// (7, 14, 'sp12_h_r_3')
// (8, 14, 'sp12_h_r_4')
// (9, 14, 'sp12_h_r_7')
// (10, 14, 'sp12_h_r_8')
// (11, 14, 'sp12_h_r_11')
// (12, 14, 'sp12_h_r_12')
// (13, 14, 'sp12_h_r_15')
// (14, 14, 'sp12_h_r_16')
// (15, 13, 'neigh_op_tnr_6')
// (15, 14, 'neigh_op_rgt_6')
// (15, 14, 'sp12_h_r_19')
// (15, 15, 'neigh_op_bnr_6')
// (16, 13, 'neigh_op_top_6')
// (16, 14, 'lutff_6/out')
// (16, 14, 'sp12_h_r_20')
// (16, 15, 'neigh_op_bot_6')
// (17, 13, 'neigh_op_tnl_6')
// (17, 14, 'neigh_op_lft_6')
// (17, 14, 'sp12_h_r_23')
// (17, 15, 'neigh_op_bnl_6')
// (18, 14, 'sp12_h_l_23')
// (18, 14, 'sp12_h_r_0')
// (19, 14, 'sp12_h_r_3')
// (20, 14, 'sp12_h_r_4')
// (21, 14, 'sp12_h_r_7')
// (22, 14, 'sp12_h_r_8')
// (23, 14, 'local_g1_3')
// (23, 14, 'lutff_global/cen')
// (23, 14, 'sp12_h_r_11')
// (24, 14, 'sp12_h_r_12')
// (25, 14, 'sp12_h_r_15')
// (26, 14, 'sp12_h_r_16')
// (27, 14, 'sp12_h_r_19')
// (28, 14, 'sp12_h_r_20')
// (29, 14, 'sp12_h_r_23')
// (30, 14, 'sp12_h_l_23')

wire n128;
// (6, 17, 'sp12_h_r_1')
// (7, 17, 'sp12_h_r_2')
// (8, 17, 'sp12_h_r_5')
// (9, 17, 'sp12_h_r_6')
// (10, 16, 'neigh_op_tnr_1')
// (10, 17, 'neigh_op_rgt_1')
// (10, 17, 'sp12_h_r_9')
// (10, 17, 'sp4_h_r_4')
// (10, 18, 'neigh_op_bnr_1')
// (11, 16, 'neigh_op_top_1')
// (11, 17, 'lutff_1/out')
// (11, 17, 'sp12_h_r_10')
// (11, 17, 'sp4_h_r_17')
// (11, 18, 'neigh_op_bot_1')
// (11, 18, 'sp4_r_v_b_37')
// (11, 19, 'sp4_r_v_b_24')
// (11, 20, 'sp4_r_v_b_13')
// (11, 21, 'sp4_r_v_b_0')
// (12, 16, 'neigh_op_tnl_1')
// (12, 17, 'local_g2_4')
// (12, 17, 'lutff_global/s_r')
// (12, 17, 'neigh_op_lft_1')
// (12, 17, 'sp12_h_r_13')
// (12, 17, 'sp4_h_r_28')
// (12, 17, 'sp4_h_r_6')
// (12, 17, 'sp4_v_t_37')
// (12, 18, 'local_g3_5')
// (12, 18, 'lutff_global/s_r')
// (12, 18, 'neigh_op_bnl_1')
// (12, 18, 'sp4_v_b_37')
// (12, 19, 'sp4_v_b_24')
// (12, 20, 'sp4_v_b_13')
// (12, 21, 'sp4_v_b_0')
// (13, 17, 'sp12_h_r_14')
// (13, 17, 'sp4_h_r_19')
// (13, 17, 'sp4_h_r_41')
// (14, 17, 'sp12_h_r_17')
// (14, 17, 'sp4_h_l_41')
// (14, 17, 'sp4_h_r_30')
// (15, 17, 'sp12_h_r_18')
// (15, 17, 'sp4_h_r_43')
// (16, 17, 'sp12_h_r_21')
// (16, 17, 'sp4_h_l_43')
// (17, 17, 'sp12_h_r_22')
// (18, 17, 'sp12_h_l_22')

reg n129 = 0;
// (6, 17, 'sp4_h_r_9')
// (7, 17, 'sp4_h_r_20')
// (8, 16, 'neigh_op_tnr_6')
// (8, 17, 'neigh_op_rgt_6')
// (8, 17, 'sp4_h_r_33')
// (8, 18, 'neigh_op_bnr_6')
// (9, 16, 'neigh_op_top_6')
// (9, 17, 'lutff_6/out')
// (9, 17, 'sp4_h_r_44')
// (9, 18, 'neigh_op_bot_6')
// (10, 16, 'neigh_op_tnl_6')
// (10, 17, 'neigh_op_lft_6')
// (10, 17, 'sp4_h_l_44')
// (10, 17, 'sp4_h_r_0')
// (10, 18, 'neigh_op_bnl_6')
// (11, 17, 'sp4_h_r_13')
// (12, 17, 'sp4_h_r_24')
// (13, 17, 'sp4_h_r_37')
// (13, 18, 'local_g2_5')
// (13, 18, 'lutff_2/in_1')
// (13, 18, 'sp4_r_v_b_37')
// (13, 19, 'sp4_r_v_b_24')
// (13, 20, 'sp4_r_v_b_13')
// (13, 21, 'sp4_r_v_b_0')
// (14, 17, 'sp4_h_l_37')
// (14, 17, 'sp4_v_t_37')
// (14, 18, 'sp4_v_b_37')
// (14, 19, 'sp4_v_b_24')
// (14, 20, 'sp4_v_b_13')
// (14, 21, 'sp4_v_b_0')

wire n130;
// (6, 18, 'sp12_h_r_1')
// (7, 18, 'sp12_h_r_2')
// (8, 18, 'sp12_h_r_5')
// (9, 18, 'sp12_h_r_6')
// (10, 18, 'sp12_h_r_9')
// (11, 18, 'sp12_h_r_10')
// (12, 17, 'neigh_op_tnr_3')
// (12, 18, 'neigh_op_rgt_3')
// (12, 18, 'sp12_h_r_13')
// (12, 19, 'neigh_op_bnr_3')
// (13, 17, 'neigh_op_top_3')
// (13, 18, 'local_g2_3')
// (13, 18, 'lutff_3/in_2')
// (13, 18, 'lutff_3/out')
// (13, 18, 'sp12_h_r_14')
// (13, 19, 'neigh_op_bot_3')
// (14, 17, 'neigh_op_tnl_3')
// (14, 18, 'neigh_op_lft_3')
// (14, 18, 'sp12_h_r_17')
// (14, 19, 'neigh_op_bnl_3')
// (15, 18, 'sp12_h_r_18')
// (16, 18, 'sp12_h_r_21')
// (17, 18, 'local_g0_6')
// (17, 18, 'lutff_3/in_1')
// (17, 18, 'sp12_h_r_22')
// (18, 18, 'sp12_h_l_22')

wire n131;
// (6, 19, 'sp12_h_r_1')
// (7, 19, 'sp12_h_r_2')
// (8, 19, 'sp12_h_r_5')
// (9, 19, 'sp12_h_r_6')
// (10, 19, 'sp12_h_r_9')
// (11, 19, 'sp12_h_r_10')
// (12, 18, 'neigh_op_tnr_3')
// (12, 19, 'neigh_op_rgt_3')
// (12, 19, 'sp12_h_r_13')
// (12, 20, 'neigh_op_bnr_3')
// (13, 18, 'neigh_op_top_3')
// (13, 19, 'local_g1_3')
// (13, 19, 'lutff_3/in_1')
// (13, 19, 'lutff_3/out')
// (13, 19, 'sp12_h_r_14')
// (13, 20, 'neigh_op_bot_3')
// (14, 18, 'neigh_op_tnl_3')
// (14, 19, 'neigh_op_lft_3')
// (14, 19, 'sp12_h_r_17')
// (14, 20, 'neigh_op_bnl_3')
// (15, 19, 'sp12_h_r_18')
// (16, 19, 'sp12_h_r_21')
// (17, 19, 'local_g0_6')
// (17, 19, 'lutff_3/in_1')
// (17, 19, 'sp12_h_r_22')
// (18, 19, 'sp12_h_l_22')

reg n132 = 0;
// (6, 24, 'sp12_h_r_0')
// (7, 24, 'sp12_h_r_3')
// (8, 24, 'sp12_h_r_4')
// (9, 24, 'sp12_h_r_7')
// (10, 24, 'sp12_h_r_8')
// (11, 24, 'sp12_h_r_11')
// (12, 24, 'sp12_h_r_12')
// (13, 24, 'sp12_h_r_15')
// (14, 24, 'sp12_h_r_16')
// (15, 23, 'neigh_op_tnr_6')
// (15, 24, 'neigh_op_rgt_6')
// (15, 24, 'sp12_h_r_19')
// (15, 25, 'neigh_op_bnr_6')
// (16, 23, 'neigh_op_top_6')
// (16, 24, 'lutff_6/out')
// (16, 24, 'sp12_h_r_20')
// (16, 25, 'neigh_op_bot_6')
// (17, 23, 'neigh_op_tnl_6')
// (17, 24, 'neigh_op_lft_6')
// (17, 24, 'sp12_h_r_23')
// (17, 25, 'neigh_op_bnl_6')
// (18, 24, 'sp12_h_l_23')
// (18, 24, 'sp12_h_r_0')
// (19, 24, 'sp12_h_r_3')
// (20, 24, 'sp12_h_r_4')
// (21, 24, 'sp12_h_r_7')
// (22, 24, 'sp12_h_r_8')
// (23, 24, 'sp12_h_r_11')
// (24, 24, 'sp12_h_r_12')
// (25, 24, 'sp12_h_r_15')
// (26, 24, 'sp12_h_r_16')
// (27, 24, 'sp12_h_r_19')
// (28, 24, 'sp12_h_r_20')
// (29, 13, 'sp4_r_v_b_45')
// (29, 14, 'sp4_r_v_b_32')
// (29, 15, 'sp4_r_v_b_21')
// (29, 16, 'sp4_r_v_b_8')
// (29, 24, 'sp12_h_r_23')
// (30, 12, 'sp12_v_t_23')
// (30, 12, 'sp4_v_t_45')
// (30, 13, 'sp12_v_b_23')
// (30, 13, 'sp4_v_b_45')
// (30, 14, 'sp12_v_b_20')
// (30, 14, 'sp4_v_b_32')
// (30, 15, 'sp12_v_b_19')
// (30, 15, 'sp4_v_b_21')
// (30, 16, 'sp12_v_b_16')
// (30, 16, 'sp4_h_r_2')
// (30, 16, 'sp4_v_b_8')
// (30, 17, 'sp12_v_b_15')
// (30, 18, 'sp12_v_b_12')
// (30, 19, 'sp12_v_b_11')
// (30, 20, 'sp12_v_b_8')
// (30, 21, 'sp12_v_b_7')
// (30, 22, 'sp12_v_b_4')
// (30, 23, 'sp12_v_b_3')
// (30, 24, 'sp12_h_l_23')
// (30, 24, 'sp12_v_b_0')
// (31, 16, 'sp4_h_r_15')
// (32, 16, 'sp4_h_r_26')
// (33, 16, 'io_1/D_OUT_0')
// (33, 16, 'local_g1_2')
// (33, 16, 'span4_horz_26')

wire io_7_33_0;
// (6, 32, 'neigh_op_tnr_0')
// (6, 32, 'neigh_op_tnr_4')
// (7, 25, 'sp12_h_r_0')
// (7, 25, 'sp12_v_t_23')
// (7, 26, 'sp12_v_b_23')
// (7, 27, 'sp12_v_b_20')
// (7, 28, 'sp12_v_b_19')
// (7, 29, 'sp12_v_b_16')
// (7, 30, 'sp12_v_b_15')
// (7, 31, 'sp12_v_b_12')
// (7, 32, 'neigh_op_top_0')
// (7, 32, 'neigh_op_top_4')
// (7, 32, 'sp12_v_b_11')
// (7, 33, 'io_0/D_IN_0')
// (7, 33, 'io_0/PAD')
// (7, 33, 'span12_vert_8')
// (8, 25, 'sp12_h_r_3')
// (8, 32, 'neigh_op_tnl_0')
// (8, 32, 'neigh_op_tnl_4')
// (9, 25, 'sp12_h_r_4')
// (10, 25, 'sp12_h_r_7')
// (11, 25, 'sp12_h_r_8')
// (12, 25, 'sp12_h_r_11')
// (12, 25, 'sp4_h_r_7')
// (13, 25, 'sp12_h_r_12')
// (13, 25, 'sp4_h_r_18')
// (14, 25, 'sp12_h_r_15')
// (14, 25, 'sp4_h_r_31')
// (15, 22, 'sp4_r_v_b_36')
// (15, 23, 'sp4_r_v_b_25')
// (15, 24, 'sp4_r_v_b_12')
// (15, 25, 'sp12_h_r_16')
// (15, 25, 'sp4_h_r_42')
// (15, 25, 'sp4_r_v_b_1')
// (16, 21, 'sp4_v_t_36')
// (16, 22, 'sp4_v_b_36')
// (16, 23, 'sp4_v_b_25')
// (16, 24, 'local_g1_4')
// (16, 24, 'lutff_0/in_3')
// (16, 24, 'sp4_v_b_12')
// (16, 25, 'sp12_h_r_19')
// (16, 25, 'sp4_h_l_42')
// (16, 25, 'sp4_v_b_1')
// (17, 25, 'sp12_h_r_20')
// (18, 25, 'sp12_h_r_23')
// (19, 25, 'sp12_h_l_23')

wire io_7_33_1;
// (6, 32, 'neigh_op_tnr_2')
// (6, 32, 'neigh_op_tnr_6')
// (7, 23, 'sp12_h_r_0')
// (7, 23, 'sp12_v_t_23')
// (7, 24, 'sp12_v_b_23')
// (7, 25, 'sp12_v_b_20')
// (7, 26, 'sp12_v_b_19')
// (7, 27, 'sp12_v_b_16')
// (7, 28, 'sp12_v_b_15')
// (7, 29, 'sp12_v_b_12')
// (7, 30, 'sp12_v_b_11')
// (7, 31, 'sp12_v_b_8')
// (7, 32, 'neigh_op_top_2')
// (7, 32, 'neigh_op_top_6')
// (7, 32, 'sp12_v_b_7')
// (7, 33, 'io_1/D_IN_0')
// (7, 33, 'io_1/PAD')
// (7, 33, 'span12_vert_4')
// (8, 23, 'sp12_h_r_3')
// (8, 32, 'neigh_op_tnl_2')
// (8, 32, 'neigh_op_tnl_6')
// (9, 23, 'sp12_h_r_4')
// (10, 23, 'sp12_h_r_7')
// (11, 23, 'sp12_h_r_8')
// (12, 23, 'sp12_h_r_11')
// (13, 23, 'sp12_h_r_12')
// (14, 23, 'sp12_h_r_15')
// (15, 23, 'sp12_h_r_16')
// (16, 23, 'local_g1_3')
// (16, 23, 'lutff_7/in_3')
// (16, 23, 'sp12_h_r_19')
// (17, 23, 'sp12_h_r_20')
// (18, 23, 'sp12_h_r_23')
// (19, 23, 'sp12_h_l_23')

reg n135 = 0;
// (7, 9, 'sp12_h_r_0')
// (8, 9, 'sp12_h_r_3')
// (9, 9, 'sp12_h_r_4')
// (10, 9, 'sp12_h_r_7')
// (11, 9, 'sp12_h_r_8')
// (12, 9, 'sp12_h_r_11')
// (13, 9, 'sp12_h_r_12')
// (14, 9, 'sp12_h_r_15')
// (15, 9, 'sp12_h_r_16')
// (16, 9, 'sp12_h_r_19')
// (17, 9, 'sp12_h_r_20')
// (18, 9, 'local_g0_7')
// (18, 9, 'lutff_0/in_3')
// (18, 9, 'sp12_h_r_23')
// (18, 20, 'neigh_op_tnr_0')
// (18, 21, 'neigh_op_rgt_0')
// (18, 22, 'neigh_op_bnr_0')
// (19, 9, 'sp12_h_l_23')
// (19, 9, 'sp12_v_t_23')
// (19, 10, 'sp12_v_b_23')
// (19, 11, 'sp12_v_b_20')
// (19, 12, 'sp12_v_b_19')
// (19, 13, 'sp12_v_b_16')
// (19, 14, 'sp12_v_b_15')
// (19, 15, 'sp12_v_b_12')
// (19, 16, 'sp12_v_b_11')
// (19, 17, 'sp12_v_b_8')
// (19, 18, 'sp12_v_b_7')
// (19, 19, 'sp12_v_b_4')
// (19, 20, 'neigh_op_top_0')
// (19, 20, 'sp12_v_b_3')
// (19, 21, 'lutff_0/out')
// (19, 21, 'sp12_v_b_0')
// (19, 22, 'neigh_op_bot_0')
// (20, 20, 'neigh_op_tnl_0')
// (20, 21, 'neigh_op_lft_0')
// (20, 22, 'neigh_op_bnl_0')

reg n136 = 0;
// (7, 10, 'local_g1_7')
// (7, 10, 'lutff_7/in_1')
// (7, 10, 'sp4_h_r_7')
// (8, 10, 'sp4_h_r_18')
// (9, 10, 'local_g3_7')
// (9, 10, 'lutff_3/in_1')
// (9, 10, 'sp4_h_r_31')
// (10, 7, 'sp4_r_v_b_42')
// (10, 8, 'neigh_op_tnr_1')
// (10, 8, 'sp4_r_v_b_31')
// (10, 9, 'local_g2_1')
// (10, 9, 'lutff_3/in_0')
// (10, 9, 'neigh_op_rgt_1')
// (10, 9, 'sp4_r_v_b_18')
// (10, 10, 'neigh_op_bnr_1')
// (10, 10, 'sp4_h_r_42')
// (10, 10, 'sp4_r_v_b_7')
// (10, 11, 'sp4_r_v_b_42')
// (10, 12, 'local_g1_7')
// (10, 12, 'lutff_1/in_1')
// (10, 12, 'sp4_r_v_b_31')
// (10, 13, 'sp4_r_v_b_18')
// (10, 14, 'sp4_r_v_b_7')
// (11, 6, 'sp4_v_t_42')
// (11, 7, 'sp4_v_b_42')
// (11, 8, 'neigh_op_top_1')
// (11, 8, 'sp4_v_b_31')
// (11, 9, 'lutff_1/out')
// (11, 9, 'sp4_v_b_18')
// (11, 10, 'neigh_op_bot_1')
// (11, 10, 'sp4_h_l_42')
// (11, 10, 'sp4_v_b_7')
// (11, 10, 'sp4_v_t_42')
// (11, 11, 'sp4_v_b_42')
// (11, 12, 'sp4_v_b_31')
// (11, 13, 'sp4_v_b_18')
// (11, 14, 'sp4_v_b_7')
// (12, 8, 'neigh_op_tnl_1')
// (12, 9, 'neigh_op_lft_1')
// (12, 10, 'neigh_op_bnl_1')

wire n137;
// (7, 12, 'lutff_6/lout')
// (7, 12, 'lutff_7/in_2')

wire n138;
// (7, 13, 'sp4_h_r_6')
// (8, 13, 'sp4_h_r_19')
// (9, 11, 'neigh_op_tnr_1')
// (9, 12, 'neigh_op_rgt_1')
// (9, 13, 'neigh_op_bnr_1')
// (9, 13, 'sp4_h_r_30')
// (10, 10, 'sp4_r_v_b_43')
// (10, 11, 'neigh_op_top_1')
// (10, 11, 'sp4_r_v_b_30')
// (10, 12, 'lutff_1/out')
// (10, 12, 'sp4_r_v_b_19')
// (10, 13, 'local_g3_3')
// (10, 13, 'lutff_global/cen')
// (10, 13, 'neigh_op_bot_1')
// (10, 13, 'sp4_h_r_43')
// (10, 13, 'sp4_r_v_b_6')
// (11, 9, 'sp4_v_t_43')
// (11, 10, 'sp4_v_b_43')
// (11, 11, 'neigh_op_tnl_1')
// (11, 11, 'sp4_v_b_30')
// (11, 12, 'neigh_op_lft_1')
// (11, 12, 'sp4_v_b_19')
// (11, 13, 'neigh_op_bnl_1')
// (11, 13, 'sp4_h_l_43')
// (11, 13, 'sp4_v_b_6')

reg n139 = 0;
// (7, 15, 'sp12_h_r_1')
// (8, 15, 'sp12_h_r_2')
// (9, 15, 'sp12_h_r_5')
// (10, 15, 'sp12_h_r_6')
// (11, 15, 'sp12_h_r_9')
// (12, 15, 'sp12_h_r_10')
// (13, 15, 'sp12_h_r_13')
// (14, 15, 'sp12_h_r_14')
// (15, 15, 'sp12_h_r_17')
// (16, 15, 'sp12_h_r_18')
// (17, 15, 'local_g1_5')
// (17, 15, 'lutff_7/in_3')
// (17, 15, 'sp12_h_r_21')
// (18, 15, 'sp12_h_r_22')
// (19, 15, 'sp12_h_l_22')
// (19, 15, 'sp12_h_r_1')
// (20, 15, 'sp12_h_r_2')
// (21, 15, 'sp12_h_r_5')
// (22, 15, 'sp12_h_r_6')
// (23, 14, 'neigh_op_tnr_1')
// (23, 15, 'neigh_op_rgt_1')
// (23, 15, 'sp12_h_r_9')
// (23, 16, 'neigh_op_bnr_1')
// (24, 14, 'neigh_op_top_1')
// (24, 15, 'lutff_1/out')
// (24, 15, 'sp12_h_r_10')
// (24, 16, 'neigh_op_bot_1')
// (25, 14, 'neigh_op_tnl_1')
// (25, 15, 'neigh_op_lft_1')
// (25, 15, 'sp12_h_r_13')
// (25, 16, 'neigh_op_bnl_1')
// (26, 15, 'sp12_h_r_14')
// (27, 15, 'sp12_h_r_17')
// (28, 15, 'sp12_h_r_18')
// (29, 15, 'sp12_h_r_21')
// (30, 15, 'sp12_h_r_22')
// (31, 15, 'sp12_h_l_22')

reg n140 = 0;
// (7, 15, 'sp4_h_r_2')
// (8, 15, 'sp4_h_r_15')
// (8, 17, 'sp4_r_v_b_41')
// (8, 18, 'sp4_r_v_b_28')
// (8, 19, 'sp4_r_v_b_17')
// (8, 20, 'sp4_r_v_b_4')
// (9, 12, 'sp12_h_r_0')
// (9, 12, 'sp12_v_t_23')
// (9, 13, 'sp12_v_b_23')
// (9, 14, 'sp12_v_b_20')
// (9, 15, 'local_g2_2')
// (9, 15, 'lutff_5/in_1')
// (9, 15, 'sp12_v_b_19')
// (9, 15, 'sp4_h_r_26')
// (9, 16, 'sp12_v_b_16')
// (9, 16, 'sp4_v_t_41')
// (9, 17, 'sp12_v_b_15')
// (9, 17, 'sp4_v_b_41')
// (9, 18, 'local_g3_4')
// (9, 18, 'lutff_2/in_3')
// (9, 18, 'sp12_v_b_12')
// (9, 18, 'sp4_v_b_28')
// (9, 19, 'sp12_v_b_11')
// (9, 19, 'sp4_v_b_17')
// (9, 20, 'sp12_v_b_8')
// (9, 20, 'sp4_h_r_10')
// (9, 20, 'sp4_v_b_4')
// (9, 21, 'sp12_v_b_7')
// (9, 22, 'sp12_v_b_4')
// (9, 23, 'sp12_v_b_3')
// (9, 24, 'sp12_v_b_0')
// (10, 11, 'neigh_op_tnr_6')
// (10, 12, 'neigh_op_rgt_6')
// (10, 12, 'sp12_h_r_3')
// (10, 12, 'sp4_h_r_1')
// (10, 12, 'sp4_r_v_b_44')
// (10, 13, 'neigh_op_bnr_6')
// (10, 13, 'sp4_r_v_b_33')
// (10, 14, 'sp4_r_v_b_20')
// (10, 15, 'sp4_h_r_39')
// (10, 15, 'sp4_r_v_b_9')
// (10, 16, 'sp4_r_v_b_44')
// (10, 17, 'sp4_r_v_b_33')
// (10, 18, 'sp4_r_v_b_20')
// (10, 19, 'local_g2_1')
// (10, 19, 'lutff_6/in_3')
// (10, 19, 'sp4_r_v_b_9')
// (10, 20, 'local_g3_0')
// (10, 20, 'lutff_4/in_3')
// (10, 20, 'sp4_h_r_23')
// (10, 20, 'sp4_r_v_b_40')
// (10, 21, 'sp4_r_v_b_29')
// (10, 22, 'sp4_r_v_b_16')
// (10, 23, 'sp4_r_v_b_5')
// (11, 10, 'sp4_r_v_b_37')
// (11, 11, 'neigh_op_top_6')
// (11, 11, 'sp4_r_v_b_24')
// (11, 11, 'sp4_v_t_44')
// (11, 12, 'lutff_6/out')
// (11, 12, 'sp12_h_r_4')
// (11, 12, 'sp4_h_r_12')
// (11, 12, 'sp4_r_v_b_13')
// (11, 12, 'sp4_v_b_44')
// (11, 13, 'local_g1_6')
// (11, 13, 'lutff_4/in_3')
// (11, 13, 'neigh_op_bot_6')
// (11, 13, 'sp4_r_v_b_0')
// (11, 13, 'sp4_v_b_33')
// (11, 14, 'sp4_v_b_20')
// (11, 15, 'sp4_h_l_39')
// (11, 15, 'sp4_v_b_9')
// (11, 15, 'sp4_v_t_44')
// (11, 16, 'sp4_v_b_44')
// (11, 17, 'sp4_v_b_33')
// (11, 18, 'sp4_v_b_20')
// (11, 19, 'sp4_h_r_9')
// (11, 19, 'sp4_v_b_9')
// (11, 19, 'sp4_v_t_40')
// (11, 20, 'sp4_h_r_34')
// (11, 20, 'sp4_v_b_40')
// (11, 21, 'sp4_v_b_29')
// (11, 22, 'local_g0_0')
// (11, 22, 'lutff_3/in_1')
// (11, 22, 'sp4_v_b_16')
// (11, 23, 'sp4_v_b_5')
// (12, 9, 'sp4_v_t_37')
// (12, 10, 'sp4_v_b_37')
// (12, 11, 'neigh_op_tnl_6')
// (12, 11, 'sp4_v_b_24')
// (12, 12, 'neigh_op_lft_6')
// (12, 12, 'sp12_h_r_7')
// (12, 12, 'sp4_h_r_25')
// (12, 12, 'sp4_v_b_13')
// (12, 13, 'local_g3_6')
// (12, 13, 'lutff_6/in_3')
// (12, 13, 'neigh_op_bnl_6')
// (12, 13, 'sp4_h_r_0')
// (12, 13, 'sp4_v_b_0')
// (12, 19, 'local_g1_4')
// (12, 19, 'lutff_6/in_3')
// (12, 19, 'sp4_h_r_20')
// (12, 20, 'local_g2_7')
// (12, 20, 'lutff_6/in_3')
// (12, 20, 'sp4_h_r_47')
// (13, 12, 'sp12_h_r_8')
// (13, 12, 'sp4_h_r_36')
// (13, 13, 'sp4_h_r_13')
// (13, 13, 'sp4_r_v_b_43')
// (13, 14, 'sp4_r_v_b_30')
// (13, 15, 'sp4_r_v_b_19')
// (13, 16, 'local_g1_6')
// (13, 16, 'lutff_4/in_3')
// (13, 16, 'sp4_r_v_b_6')
// (13, 19, 'sp4_h_r_33')
// (13, 20, 'sp4_h_l_47')
// (14, 12, 'sp12_h_r_11')
// (14, 12, 'sp4_h_l_36')
// (14, 12, 'sp4_h_r_9')
// (14, 12, 'sp4_v_t_43')
// (14, 13, 'local_g3_0')
// (14, 13, 'lutff_6/in_3')
// (14, 13, 'sp4_h_r_24')
// (14, 13, 'sp4_v_b_43')
// (14, 14, 'sp4_v_b_30')
// (14, 15, 'local_g0_3')
// (14, 15, 'lutff_1/in_0')
// (14, 15, 'sp4_v_b_19')
// (14, 16, 'sp4_v_b_6')
// (14, 19, 'sp4_h_r_44')
// (14, 20, 'sp4_r_v_b_44')
// (14, 21, 'sp4_r_v_b_33')
// (14, 22, 'local_g3_4')
// (14, 22, 'lutff_4/in_3')
// (14, 22, 'sp4_r_v_b_20')
// (14, 23, 'sp4_r_v_b_9')
// (15, 10, 'sp4_r_v_b_43')
// (15, 11, 'sp4_r_v_b_30')
// (15, 12, 'sp12_h_r_12')
// (15, 12, 'sp4_h_r_20')
// (15, 12, 'sp4_r_v_b_19')
// (15, 13, 'local_g3_5')
// (15, 13, 'lutff_7/in_3')
// (15, 13, 'sp4_h_r_37')
// (15, 13, 'sp4_r_v_b_6')
// (15, 14, 'sp4_r_v_b_37')
// (15, 15, 'local_g1_0')
// (15, 15, 'lutff_6/in_3')
// (15, 15, 'sp4_r_v_b_24')
// (15, 16, 'sp4_r_v_b_13')
// (15, 17, 'local_g1_0')
// (15, 17, 'lutff_6/in_3')
// (15, 17, 'sp4_r_v_b_0')
// (15, 18, 'local_g2_5')
// (15, 18, 'lutff_6/in_3')
// (15, 18, 'sp4_r_v_b_37')
// (15, 19, 'local_g1_0')
// (15, 19, 'lutff_6/in_3')
// (15, 19, 'sp4_h_l_44')
// (15, 19, 'sp4_r_v_b_24')
// (15, 19, 'sp4_v_t_44')
// (15, 20, 'sp4_r_v_b_13')
// (15, 20, 'sp4_v_b_44')
// (15, 21, 'sp4_r_v_b_0')
// (15, 21, 'sp4_v_b_33')
// (15, 22, 'sp4_v_b_20')
// (15, 23, 'sp4_v_b_9')
// (16, 9, 'sp4_v_t_43')
// (16, 10, 'sp4_v_b_43')
// (16, 11, 'local_g3_6')
// (16, 11, 'lutff_6/in_3')
// (16, 11, 'sp4_v_b_30')
// (16, 12, 'sp12_h_r_15')
// (16, 12, 'sp4_h_r_33')
// (16, 12, 'sp4_v_b_19')
// (16, 13, 'sp4_h_l_37')
// (16, 13, 'sp4_h_r_3')
// (16, 13, 'sp4_v_b_6')
// (16, 13, 'sp4_v_t_37')
// (16, 14, 'sp4_v_b_37')
// (16, 15, 'sp4_v_b_24')
// (16, 16, 'local_g0_5')
// (16, 16, 'lutff_6/in_3')
// (16, 16, 'sp4_v_b_13')
// (16, 17, 'local_g1_0')
// (16, 17, 'lutff_6/in_3')
// (16, 17, 'sp4_v_b_0')
// (16, 17, 'sp4_v_t_37')
// (16, 18, 'local_g2_5')
// (16, 18, 'lutff_6/in_3')
// (16, 18, 'sp4_v_b_37')
// (16, 19, 'local_g3_0')
// (16, 19, 'lutff_4/in_3')
// (16, 19, 'sp4_v_b_24')
// (16, 20, 'sp4_v_b_13')
// (16, 21, 'local_g0_0')
// (16, 21, 'lutff_4/in_0')
// (16, 21, 'sp4_v_b_0')
// (17, 9, 'sp4_r_v_b_44')
// (17, 10, 'sp4_r_v_b_33')
// (17, 11, 'local_g3_4')
// (17, 11, 'lutff_7/in_0')
// (17, 11, 'sp4_r_v_b_20')
// (17, 12, 'local_g3_4')
// (17, 12, 'lutff_0/in_3')
// (17, 12, 'sp12_h_r_16')
// (17, 12, 'sp4_h_r_44')
// (17, 12, 'sp4_r_v_b_9')
// (17, 13, 'local_g1_6')
// (17, 13, 'lutff_0/in_3')
// (17, 13, 'sp4_h_r_14')
// (17, 13, 'sp4_r_v_b_39')
// (17, 14, 'local_g1_2')
// (17, 14, 'lutff_5/in_0')
// (17, 14, 'sp4_r_v_b_26')
// (17, 15, 'local_g2_7')
// (17, 15, 'lutff_2/in_3')
// (17, 15, 'sp4_r_v_b_15')
// (17, 16, 'sp4_r_v_b_2')
// (17, 17, 'sp4_r_v_b_39')
// (17, 18, 'sp4_r_v_b_26')
// (17, 19, 'sp4_r_v_b_15')
// (17, 20, 'sp4_r_v_b_2')
// (18, 8, 'sp4_v_t_44')
// (18, 9, 'sp4_v_b_44')
// (18, 10, 'sp4_v_b_33')
// (18, 11, 'sp4_v_b_20')
// (18, 12, 'local_g0_3')
// (18, 12, 'lutff_6/in_3')
// (18, 12, 'sp12_h_r_19')
// (18, 12, 'sp4_h_l_44')
// (18, 12, 'sp4_v_b_9')
// (18, 12, 'sp4_v_t_39')
// (18, 13, 'sp4_h_r_27')
// (18, 13, 'sp4_v_b_39')
// (18, 14, 'sp4_v_b_26')
// (18, 15, 'sp4_v_b_15')
// (18, 16, 'sp4_h_r_8')
// (18, 16, 'sp4_v_b_2')
// (18, 16, 'sp4_v_t_39')
// (18, 17, 'sp4_v_b_39')
// (18, 18, 'sp4_v_b_26')
// (18, 19, 'local_g1_7')
// (18, 19, 'lutff_1/in_3')
// (18, 19, 'sp4_v_b_15')
// (18, 20, 'sp4_h_r_8')
// (18, 20, 'sp4_v_b_2')
// (19, 10, 'local_g3_4')
// (19, 10, 'lutff_6/in_3')
// (19, 10, 'sp4_r_v_b_44')
// (19, 11, 'local_g2_1')
// (19, 11, 'lutff_6/in_3')
// (19, 11, 'sp4_r_v_b_33')
// (19, 12, 'sp12_h_r_20')
// (19, 12, 'sp4_r_v_b_20')
// (19, 13, 'sp4_h_r_38')
// (19, 13, 'sp4_r_v_b_9')
// (19, 14, 'sp4_r_v_b_38')
// (19, 15, 'sp4_r_v_b_27')
// (19, 16, 'local_g0_5')
// (19, 16, 'lutff_6/in_3')
// (19, 16, 'sp4_h_r_21')
// (19, 16, 'sp4_r_v_b_14')
// (19, 17, 'sp4_r_v_b_3')
// (19, 18, 'sp4_r_v_b_46')
// (19, 19, 'local_g0_0')
// (19, 19, 'lutff_5/in_1')
// (19, 19, 'sp4_r_v_b_35')
// (19, 20, 'sp4_h_r_21')
// (19, 20, 'sp4_r_v_b_22')
// (19, 21, 'sp4_r_v_b_11')
// (19, 22, 'sp4_r_v_b_46')
// (19, 23, 'sp4_r_v_b_35')
// (19, 24, 'sp4_r_v_b_22')
// (19, 25, 'sp4_r_v_b_11')
// (20, 9, 'sp4_v_t_44')
// (20, 10, 'sp4_v_b_44')
// (20, 11, 'local_g3_1')
// (20, 11, 'lutff_5/in_3')
// (20, 11, 'sp4_v_b_33')
// (20, 12, 'local_g0_7')
// (20, 12, 'lutff_6/in_3')
// (20, 12, 'sp12_h_r_23')
// (20, 12, 'sp4_v_b_20')
// (20, 13, 'sp4_h_l_38')
// (20, 13, 'sp4_h_r_3')
// (20, 13, 'sp4_v_b_9')
// (20, 13, 'sp4_v_t_38')
// (20, 14, 'sp4_v_b_38')
// (20, 15, 'sp4_v_b_27')
// (20, 16, 'local_g3_0')
// (20, 16, 'lutff_6/in_3')
// (20, 16, 'sp4_h_r_32')
// (20, 16, 'sp4_v_b_14')
// (20, 17, 'sp4_v_b_3')
// (20, 17, 'sp4_v_t_46')
// (20, 18, 'sp4_v_b_46')
// (20, 19, 'local_g2_3')
// (20, 19, 'lutff_6/in_3')
// (20, 19, 'sp4_v_b_35')
// (20, 20, 'local_g1_6')
// (20, 20, 'lutff_6/in_3')
// (20, 20, 'sp4_h_r_32')
// (20, 20, 'sp4_v_b_22')
// (20, 21, 'local_g1_5')
// (20, 21, 'lutff_7/in_3')
// (20, 21, 'sp4_h_r_5')
// (20, 21, 'sp4_v_b_11')
// (20, 21, 'sp4_v_t_46')
// (20, 22, 'sp4_v_b_46')
// (20, 23, 'sp4_v_b_35')
// (20, 24, 'sp4_v_b_22')
// (20, 25, 'local_g0_3')
// (20, 25, 'lutff_6/in_3')
// (20, 25, 'sp4_v_b_11')
// (21, 0, 'span12_vert_23')
// (21, 1, 'sp12_v_b_23')
// (21, 2, 'sp12_v_b_20')
// (21, 3, 'sp12_v_b_19')
// (21, 4, 'sp12_v_b_16')
// (21, 5, 'sp12_v_b_15')
// (21, 6, 'sp12_v_b_12')
// (21, 7, 'sp12_v_b_11')
// (21, 8, 'sp12_v_b_8')
// (21, 9, 'sp12_v_b_7')
// (21, 10, 'sp12_v_b_4')
// (21, 11, 'local_g2_3')
// (21, 11, 'lutff_6/in_3')
// (21, 11, 'sp12_v_b_3')
// (21, 12, 'local_g1_0')
// (21, 12, 'lutff_6/in_3')
// (21, 12, 'sp12_h_l_23')
// (21, 12, 'sp12_h_r_0')
// (21, 12, 'sp12_v_b_0')
// (21, 13, 'sp4_h_r_14')
// (21, 13, 'sp4_r_v_b_45')
// (21, 14, 'sp4_r_v_b_32')
// (21, 15, 'sp4_r_v_b_21')
// (21, 16, 'sp4_h_r_45')
// (21, 16, 'sp4_r_v_b_8')
// (21, 17, 'local_g3_1')
// (21, 17, 'lutff_7/in_3')
// (21, 17, 'sp4_r_v_b_41')
// (21, 18, 'sp4_r_v_b_28')
// (21, 19, 'sp4_r_v_b_17')
// (21, 20, 'local_g2_5')
// (21, 20, 'lutff_6/in_3')
// (21, 20, 'sp4_h_r_45')
// (21, 20, 'sp4_r_v_b_4')
// (21, 21, 'sp4_h_r_16')
// (21, 21, 'sp4_r_v_b_42')
// (21, 22, 'sp4_r_v_b_31')
// (21, 23, 'sp4_r_v_b_18')
// (21, 24, 'sp4_r_v_b_7')
// (22, 12, 'local_g0_3')
// (22, 12, 'lutff_6/in_3')
// (22, 12, 'sp12_h_r_3')
// (22, 12, 'sp4_v_t_45')
// (22, 13, 'sp4_h_r_27')
// (22, 13, 'sp4_v_b_45')
// (22, 14, 'local_g3_0')
// (22, 14, 'lutff_6/in_3')
// (22, 14, 'sp4_v_b_32')
// (22, 15, 'sp4_v_b_21')
// (22, 16, 'sp4_h_l_45')
// (22, 16, 'sp4_v_b_8')
// (22, 16, 'sp4_v_t_41')
// (22, 17, 'sp4_v_b_41')
// (22, 18, 'sp4_v_b_28')
// (22, 19, 'local_g1_1')
// (22, 19, 'lutff_5/in_3')
// (22, 19, 'sp4_v_b_17')
// (22, 20, 'sp4_h_l_45')
// (22, 20, 'sp4_v_b_4')
// (22, 20, 'sp4_v_t_42')
// (22, 21, 'local_g2_5')
// (22, 21, 'lutff_6/in_3')
// (22, 21, 'sp4_h_r_29')
// (22, 21, 'sp4_v_b_42')
// (22, 22, 'sp4_v_b_31')
// (22, 23, 'local_g1_2')
// (22, 23, 'lutff_6/in_3')
// (22, 23, 'sp4_v_b_18')
// (22, 24, 'sp4_v_b_7')
// (23, 12, 'local_g1_4')
// (23, 12, 'lutff_6/in_3')
// (23, 12, 'sp12_h_r_4')
// (23, 13, 'local_g2_6')
// (23, 13, 'lutff_5/in_3')
// (23, 13, 'sp4_h_r_38')
// (23, 14, 'local_g2_6')
// (23, 14, 'lutff_6/in_0')
// (23, 14, 'sp4_r_v_b_38')
// (23, 15, 'local_g0_3')
// (23, 15, 'lutff_6/in_3')
// (23, 15, 'sp4_r_v_b_27')
// (23, 16, 'local_g2_6')
// (23, 16, 'lutff_6/in_0')
// (23, 16, 'sp4_r_v_b_14')
// (23, 17, 'sp4_r_v_b_3')
// (23, 18, 'sp4_r_v_b_46')
// (23, 19, 'sp4_r_v_b_35')
// (23, 20, 'local_g3_6')
// (23, 20, 'lutff_6/in_3')
// (23, 20, 'sp4_r_v_b_22')
// (23, 21, 'sp4_h_r_40')
// (23, 21, 'sp4_r_v_b_11')
// (24, 12, 'sp12_h_r_7')
// (24, 13, 'sp4_h_l_38')
// (24, 13, 'sp4_v_t_38')
// (24, 14, 'local_g3_6')
// (24, 14, 'lutff_6/in_3')
// (24, 14, 'sp4_v_b_38')
// (24, 15, 'sp4_v_b_27')
// (24, 16, 'sp4_v_b_14')
// (24, 17, 'local_g1_3')
// (24, 17, 'lutff_6/in_0')
// (24, 17, 'sp4_v_b_3')
// (24, 17, 'sp4_v_t_46')
// (24, 18, 'sp4_v_b_46')
// (24, 19, 'sp4_v_b_35')
// (24, 20, 'sp4_v_b_22')
// (24, 21, 'sp4_h_l_40')
// (24, 21, 'sp4_v_b_11')
// (25, 12, 'sp12_h_r_8')
// (26, 12, 'sp12_h_r_11')
// (27, 12, 'sp12_h_r_12')
// (28, 12, 'sp12_h_r_15')
// (29, 12, 'sp12_h_r_16')
// (30, 12, 'sp12_h_r_19')
// (31, 12, 'sp12_h_r_20')
// (32, 12, 'sp12_h_r_23')
// (33, 12, 'span12_horz_23')

wire n141;
// (7, 17, 'sp4_h_r_9')
// (8, 17, 'sp4_h_r_20')
// (9, 17, 'local_g2_1')
// (9, 17, 'lutff_0/in_3')
// (9, 17, 'sp4_h_r_33')
// (10, 17, 'sp4_h_r_44')
// (11, 17, 'sp4_h_l_44')
// (11, 17, 'sp4_h_r_1')
// (12, 17, 'sp4_h_r_12')
// (13, 17, 'sp4_h_r_25')
// (14, 14, 'sp4_r_v_b_36')
// (14, 15, 'neigh_op_tnr_6')
// (14, 15, 'sp4_r_v_b_25')
// (14, 16, 'neigh_op_rgt_6')
// (14, 16, 'sp4_r_v_b_12')
// (14, 17, 'neigh_op_bnr_6')
// (14, 17, 'sp4_h_r_36')
// (14, 17, 'sp4_r_v_b_1')
// (15, 13, 'sp4_v_t_36')
// (15, 14, 'sp4_v_b_36')
// (15, 15, 'neigh_op_top_6')
// (15, 15, 'sp4_v_b_25')
// (15, 16, 'local_g2_6')
// (15, 16, 'lutff_4/in_0')
// (15, 16, 'lutff_5/in_3')
// (15, 16, 'lutff_6/out')
// (15, 16, 'sp4_v_b_12')
// (15, 17, 'neigh_op_bot_6')
// (15, 17, 'sp4_h_l_36')
// (15, 17, 'sp4_v_b_1')
// (16, 15, 'neigh_op_tnl_6')
// (16, 16, 'neigh_op_lft_6')
// (16, 17, 'neigh_op_bnl_6')

wire n142;
// (7, 18, 'sp12_h_r_0')
// (8, 18, 'sp12_h_r_3')
// (9, 18, 'sp12_h_r_4')
// (10, 18, 'sp12_h_r_7')
// (11, 18, 'sp12_h_r_8')
// (12, 17, 'neigh_op_tnr_2')
// (12, 18, 'neigh_op_rgt_2')
// (12, 18, 'sp12_h_r_11')
// (12, 19, 'neigh_op_bnr_2')
// (13, 17, 'neigh_op_top_2')
// (13, 18, 'local_g2_2')
// (13, 18, 'lutff_2/in_2')
// (13, 18, 'lutff_2/out')
// (13, 18, 'sp12_h_r_12')
// (13, 19, 'neigh_op_bot_2')
// (14, 17, 'neigh_op_tnl_2')
// (14, 18, 'neigh_op_lft_2')
// (14, 18, 'sp12_h_r_15')
// (14, 19, 'neigh_op_bnl_2')
// (15, 18, 'sp12_h_r_16')
// (16, 18, 'sp12_h_r_19')
// (17, 18, 'local_g1_4')
// (17, 18, 'lutff_2/in_1')
// (17, 18, 'sp12_h_r_20')
// (18, 18, 'sp12_h_r_23')
// (19, 18, 'sp12_h_l_23')

wire n143;
// (7, 19, 'sp12_h_r_0')
// (8, 19, 'sp12_h_r_3')
// (9, 19, 'sp12_h_r_4')
// (10, 19, 'sp12_h_r_7')
// (11, 19, 'sp12_h_r_8')
// (12, 18, 'neigh_op_tnr_2')
// (12, 19, 'neigh_op_rgt_2')
// (12, 19, 'sp12_h_r_11')
// (12, 20, 'neigh_op_bnr_2')
// (13, 18, 'neigh_op_top_2')
// (13, 19, 'local_g2_2')
// (13, 19, 'lutff_2/in_2')
// (13, 19, 'lutff_2/out')
// (13, 19, 'sp12_h_r_12')
// (13, 20, 'neigh_op_bot_2')
// (14, 18, 'neigh_op_tnl_2')
// (14, 19, 'neigh_op_lft_2')
// (14, 19, 'sp12_h_r_15')
// (14, 20, 'neigh_op_bnl_2')
// (15, 19, 'sp12_h_r_16')
// (16, 19, 'sp12_h_r_19')
// (17, 19, 'local_g1_4')
// (17, 19, 'lutff_2/in_1')
// (17, 19, 'sp12_h_r_20')
// (18, 19, 'sp12_h_r_23')
// (19, 19, 'sp12_h_l_23')

wire n144;
// (7, 20, 'sp4_h_r_7')
// (8, 20, 'sp4_h_r_18')
// (9, 20, 'sp4_h_r_31')
// (10, 20, 'local_g2_2')
// (10, 20, 'lutff_global/cen')
// (10, 20, 'sp4_h_r_42')
// (11, 20, 'sp4_h_l_42')
// (11, 20, 'sp4_h_r_4')
// (12, 20, 'sp4_h_r_17')
// (13, 20, 'sp4_h_r_28')
// (14, 20, 'sp4_h_r_41')
// (15, 19, 'neigh_op_tnr_6')
// (15, 20, 'neigh_op_rgt_6')
// (15, 20, 'sp4_h_l_41')
// (15, 20, 'sp4_h_r_1')
// (15, 21, 'neigh_op_bnr_6')
// (16, 19, 'neigh_op_top_6')
// (16, 20, 'lutff_6/out')
// (16, 20, 'sp4_h_r_12')
// (16, 21, 'neigh_op_bot_6')
// (17, 19, 'neigh_op_tnl_6')
// (17, 20, 'neigh_op_lft_6')
// (17, 20, 'sp4_h_r_25')
// (17, 21, 'neigh_op_bnl_6')
// (18, 20, 'sp4_h_r_36')
// (19, 20, 'sp4_h_l_36')

reg n145 = 0;
// (7, 22, 'sp12_h_r_0')
// (8, 22, 'sp12_h_r_3')
// (9, 22, 'sp12_h_r_4')
// (10, 21, 'neigh_op_tnr_0')
// (10, 22, 'neigh_op_rgt_0')
// (10, 22, 'sp12_h_r_7')
// (10, 23, 'neigh_op_bnr_0')
// (11, 21, 'neigh_op_top_0')
// (11, 22, 'lutff_0/out')
// (11, 22, 'sp12_h_r_8')
// (11, 23, 'neigh_op_bot_0')
// (12, 21, 'neigh_op_tnl_0')
// (12, 22, 'neigh_op_lft_0')
// (12, 22, 'sp12_h_r_11')
// (12, 23, 'neigh_op_bnl_0')
// (13, 22, 'local_g0_4')
// (13, 22, 'lutff_0/in_0')
// (13, 22, 'sp12_h_r_12')
// (14, 22, 'sp12_h_r_15')
// (15, 22, 'sp12_h_r_16')
// (16, 22, 'sp12_h_r_19')
// (17, 22, 'sp12_h_r_20')
// (18, 22, 'sp12_h_r_23')
// (19, 22, 'sp12_h_l_23')

reg n146 = 0;
// (7, 24, 'sp12_h_r_1')
// (8, 24, 'sp12_h_r_2')
// (9, 24, 'sp12_h_r_5')
// (10, 24, 'sp12_h_r_6')
// (11, 24, 'sp12_h_r_9')
// (12, 24, 'sp12_h_r_10')
// (13, 24, 'sp12_h_r_13')
// (14, 24, 'sp12_h_r_14')
// (15, 23, 'neigh_op_tnr_5')
// (15, 24, 'neigh_op_rgt_5')
// (15, 24, 'sp12_h_r_17')
// (15, 25, 'neigh_op_bnr_5')
// (16, 23, 'neigh_op_top_5')
// (16, 24, 'lutff_5/out')
// (16, 24, 'sp12_h_r_18')
// (16, 25, 'neigh_op_bot_5')
// (17, 23, 'neigh_op_tnl_5')
// (17, 24, 'neigh_op_lft_5')
// (17, 24, 'sp12_h_r_21')
// (17, 25, 'neigh_op_bnl_5')
// (18, 24, 'sp12_h_r_22')
// (19, 24, 'sp12_h_l_22')
// (19, 24, 'sp12_h_r_1')
// (20, 24, 'sp12_h_r_2')
// (21, 24, 'sp12_h_r_5')
// (22, 24, 'sp12_h_r_6')
// (23, 24, 'sp12_h_r_9')
// (24, 24, 'sp12_h_r_10')
// (25, 24, 'sp12_h_r_13')
// (26, 24, 'sp12_h_r_14')
// (27, 24, 'sp12_h_r_17')
// (28, 24, 'sp12_h_r_18')
// (29, 24, 'sp12_h_r_21')
// (30, 24, 'sp12_h_r_22')
// (31, 12, 'sp12_h_r_1')
// (31, 12, 'sp12_v_t_22')
// (31, 12, 'sp4_h_r_0')
// (31, 13, 'sp12_v_b_22')
// (31, 14, 'sp12_v_b_21')
// (31, 15, 'sp12_v_b_18')
// (31, 16, 'sp12_v_b_17')
// (31, 17, 'sp12_v_b_14')
// (31, 18, 'sp12_v_b_13')
// (31, 19, 'sp12_v_b_10')
// (31, 20, 'sp12_v_b_9')
// (31, 21, 'sp12_v_b_6')
// (31, 22, 'sp12_v_b_5')
// (31, 23, 'sp12_v_b_2')
// (31, 24, 'sp12_h_l_22')
// (31, 24, 'sp12_v_b_1')
// (32, 12, 'sp12_h_r_2')
// (32, 12, 'sp4_h_r_13')
// (33, 8, 'span4_vert_t_14')
// (33, 9, 'span4_vert_b_14')
// (33, 10, 'io_1/D_OUT_0')
// (33, 10, 'local_g1_2')
// (33, 10, 'span4_vert_b_10')
// (33, 11, 'span4_vert_b_6')
// (33, 12, 'span12_horz_2')
// (33, 12, 'span4_horz_13')
// (33, 12, 'span4_vert_b_2')

wire io_8_33_0;
// (7, 32, 'neigh_op_tnr_0')
// (7, 32, 'neigh_op_tnr_4')
// (8, 25, 'sp12_h_r_0')
// (8, 25, 'sp12_v_t_23')
// (8, 26, 'sp12_v_b_23')
// (8, 27, 'sp12_v_b_20')
// (8, 28, 'sp12_v_b_19')
// (8, 29, 'sp12_v_b_16')
// (8, 30, 'sp12_v_b_15')
// (8, 31, 'sp12_v_b_12')
// (8, 32, 'neigh_op_top_0')
// (8, 32, 'neigh_op_top_4')
// (8, 32, 'sp12_v_b_11')
// (8, 33, 'io_0/D_IN_0')
// (8, 33, 'io_0/PAD')
// (8, 33, 'span12_vert_8')
// (9, 25, 'sp12_h_r_3')
// (9, 32, 'neigh_op_tnl_0')
// (9, 32, 'neigh_op_tnl_4')
// (10, 25, 'sp12_h_r_4')
// (11, 25, 'sp12_h_r_7')
// (12, 25, 'sp12_h_r_8')
// (13, 25, 'sp12_h_r_11')
// (13, 25, 'sp4_h_r_7')
// (14, 25, 'sp12_h_r_12')
// (14, 25, 'sp4_h_r_18')
// (15, 25, 'sp12_h_r_15')
// (15, 25, 'sp4_h_r_31')
// (16, 22, 'sp4_r_v_b_42')
// (16, 23, 'local_g1_7')
// (16, 23, 'lutff_1/in_3')
// (16, 23, 'sp4_r_v_b_31')
// (16, 24, 'sp4_r_v_b_18')
// (16, 25, 'sp12_h_r_16')
// (16, 25, 'sp4_h_r_42')
// (16, 25, 'sp4_r_v_b_7')
// (17, 21, 'sp4_v_t_42')
// (17, 22, 'sp4_v_b_42')
// (17, 23, 'sp4_v_b_31')
// (17, 24, 'sp4_v_b_18')
// (17, 25, 'sp12_h_r_19')
// (17, 25, 'sp4_h_l_42')
// (17, 25, 'sp4_v_b_7')
// (18, 25, 'sp12_h_r_20')
// (19, 25, 'sp12_h_r_23')
// (20, 25, 'sp12_h_l_23')

wire io_8_33_1;
// (7, 32, 'neigh_op_tnr_2')
// (7, 32, 'neigh_op_tnr_6')
// (8, 23, 'sp12_h_r_0')
// (8, 23, 'sp12_v_t_23')
// (8, 24, 'sp12_v_b_23')
// (8, 25, 'sp12_v_b_20')
// (8, 26, 'sp12_v_b_19')
// (8, 27, 'sp12_v_b_16')
// (8, 28, 'sp12_v_b_15')
// (8, 29, 'sp12_v_b_12')
// (8, 30, 'sp12_v_b_11')
// (8, 31, 'sp12_v_b_8')
// (8, 32, 'neigh_op_top_2')
// (8, 32, 'neigh_op_top_6')
// (8, 32, 'sp12_v_b_7')
// (8, 33, 'io_1/D_IN_0')
// (8, 33, 'io_1/PAD')
// (8, 33, 'span12_vert_4')
// (9, 23, 'sp12_h_r_3')
// (9, 32, 'neigh_op_tnl_2')
// (9, 32, 'neigh_op_tnl_6')
// (10, 23, 'sp12_h_r_4')
// (11, 23, 'sp12_h_r_7')
// (12, 23, 'sp12_h_r_8')
// (13, 23, 'sp12_h_r_11')
// (14, 23, 'sp12_h_r_12')
// (15, 23, 'sp12_h_r_15')
// (16, 23, 'local_g1_0')
// (16, 23, 'lutff_0/in_3')
// (16, 23, 'sp12_h_r_16')
// (17, 23, 'sp12_h_r_19')
// (18, 23, 'sp12_h_r_20')
// (19, 23, 'sp12_h_r_23')
// (20, 23, 'sp12_h_l_23')

reg n149 = 0;
// (8, 8, 'sp12_h_r_1')
// (9, 8, 'sp12_h_r_2')
// (10, 8, 'sp12_h_r_5')
// (11, 8, 'sp12_h_r_6')
// (12, 8, 'sp12_h_r_9')
// (13, 8, 'local_g1_2')
// (13, 8, 'lutff_6/in_3')
// (13, 8, 'sp12_h_r_10')
// (14, 8, 'sp12_h_r_13')
// (15, 8, 'sp12_h_r_14')
// (16, 7, 'neigh_op_tnr_5')
// (16, 8, 'neigh_op_rgt_5')
// (16, 8, 'sp12_h_r_17')
// (16, 9, 'neigh_op_bnr_5')
// (17, 7, 'neigh_op_top_5')
// (17, 8, 'lutff_5/out')
// (17, 8, 'sp12_h_r_18')
// (17, 9, 'neigh_op_bot_5')
// (18, 7, 'neigh_op_tnl_5')
// (18, 8, 'neigh_op_lft_5')
// (18, 8, 'sp12_h_r_21')
// (18, 9, 'neigh_op_bnl_5')
// (19, 8, 'sp12_h_r_22')
// (20, 8, 'sp12_h_l_22')

wire n150;
// (8, 9, 'neigh_op_tnr_3')
// (8, 10, 'neigh_op_rgt_3')
// (8, 10, 'sp4_r_v_b_38')
// (8, 11, 'neigh_op_bnr_3')
// (8, 11, 'sp4_r_v_b_27')
// (8, 12, 'sp4_r_v_b_14')
// (8, 13, 'sp4_r_v_b_3')
// (9, 9, 'neigh_op_top_3')
// (9, 9, 'sp4_h_r_3')
// (9, 9, 'sp4_v_t_38')
// (9, 10, 'lutff_3/out')
// (9, 10, 'sp4_v_b_38')
// (9, 11, 'neigh_op_bot_3')
// (9, 11, 'sp4_v_b_27')
// (9, 12, 'sp4_v_b_14')
// (9, 13, 'sp4_v_b_3')
// (10, 9, 'local_g3_3')
// (10, 9, 'lutff_0/in_2')
// (10, 9, 'lutff_1/in_3')
// (10, 9, 'lutff_5/in_1')
// (10, 9, 'neigh_op_tnl_3')
// (10, 9, 'sp4_h_r_14')
// (10, 10, 'local_g1_3')
// (10, 10, 'lutff_4/in_0')
// (10, 10, 'neigh_op_lft_3')
// (10, 11, 'local_g3_3')
// (10, 11, 'lutff_global/cen')
// (10, 11, 'neigh_op_bnl_3')
// (11, 9, 'local_g2_3')
// (11, 9, 'local_g3_3')
// (11, 9, 'lutff_5/in_1')
// (11, 9, 'lutff_7/in_0')
// (11, 9, 'sp4_h_r_27')
// (12, 9, 'sp4_h_r_38')
// (13, 9, 'sp4_h_l_38')

reg n151 = 0;
// (8, 9, 'sp12_h_r_1')
// (9, 9, 'sp12_h_r_2')
// (10, 8, 'neigh_op_tnr_7')
// (10, 9, 'neigh_op_rgt_7')
// (10, 9, 'sp12_h_r_5')
// (10, 9, 'sp4_h_r_2')
// (10, 10, 'local_g0_7')
// (10, 10, 'lutff_2/in_1')
// (10, 10, 'neigh_op_bnr_7')
// (11, 8, 'neigh_op_top_7')
// (11, 9, 'local_g3_7')
// (11, 9, 'lutff_4/in_0')
// (11, 9, 'lutff_6/in_0')
// (11, 9, 'lutff_7/in_1')
// (11, 9, 'lutff_7/out')
// (11, 9, 'sp12_h_r_6')
// (11, 9, 'sp4_h_r_15')
// (11, 10, 'neigh_op_bot_7')
// (12, 8, 'neigh_op_tnl_7')
// (12, 9, 'neigh_op_lft_7')
// (12, 9, 'sp12_h_r_9')
// (12, 9, 'sp4_h_r_26')
// (12, 10, 'local_g2_7')
// (12, 10, 'lutff_2/in_3')
// (12, 10, 'neigh_op_bnl_7')
// (13, 9, 'sp12_h_r_10')
// (13, 9, 'sp4_h_r_39')
// (13, 10, 'sp4_r_v_b_42')
// (13, 11, 'sp4_r_v_b_31')
// (13, 12, 'sp4_r_v_b_18')
// (13, 13, 'sp4_r_v_b_7')
// (14, 9, 'local_g1_5')
// (14, 9, 'lutff_4/in_0')
// (14, 9, 'sp12_h_r_13')
// (14, 9, 'sp4_h_l_39')
// (14, 9, 'sp4_v_t_42')
// (14, 10, 'sp4_v_b_42')
// (14, 11, 'sp4_v_b_31')
// (14, 12, 'local_g1_2')
// (14, 12, 'lutff_1/in_0')
// (14, 12, 'lutff_3/in_0')
// (14, 12, 'sp4_v_b_18')
// (14, 13, 'sp4_v_b_7')
// (15, 9, 'sp12_h_r_14')
// (16, 9, 'sp12_h_r_17')
// (17, 9, 'sp12_h_r_18')
// (18, 9, 'sp12_h_r_21')
// (19, 9, 'sp12_h_r_22')
// (20, 9, 'sp12_h_l_22')

reg n152 = 0;
// (8, 9, 'sp4_h_r_2')
// (9, 8, 'neigh_op_tnr_5')
// (9, 9, 'neigh_op_rgt_5')
// (9, 9, 'sp12_h_r_1')
// (9, 9, 'sp4_h_r_15')
// (9, 10, 'neigh_op_bnr_5')
// (10, 8, 'neigh_op_top_5')
// (10, 9, 'local_g0_5')
// (10, 9, 'lutff_5/in_2')
// (10, 9, 'lutff_5/out')
// (10, 9, 'sp12_h_r_2')
// (10, 9, 'sp4_h_r_26')
// (10, 9, 'sp4_r_v_b_43')
// (10, 10, 'local_g1_5')
// (10, 10, 'lutff_3/in_1')
// (10, 10, 'neigh_op_bot_5')
// (10, 10, 'sp4_r_v_b_30')
// (10, 11, 'sp4_r_v_b_19')
// (10, 12, 'sp4_r_v_b_6')
// (11, 8, 'neigh_op_tnl_5')
// (11, 8, 'sp4_v_t_43')
// (11, 9, 'local_g0_5')
// (11, 9, 'lutff_4/in_1')
// (11, 9, 'lutff_6/in_3')
// (11, 9, 'neigh_op_lft_5')
// (11, 9, 'sp12_h_r_5')
// (11, 9, 'sp4_h_r_2')
// (11, 9, 'sp4_h_r_39')
// (11, 9, 'sp4_v_b_43')
// (11, 10, 'neigh_op_bnl_5')
// (11, 10, 'sp4_r_v_b_42')
// (11, 10, 'sp4_v_b_30')
// (11, 11, 'sp4_r_v_b_31')
// (11, 11, 'sp4_v_b_19')
// (11, 12, 'sp4_h_r_6')
// (11, 12, 'sp4_r_v_b_18')
// (11, 12, 'sp4_v_b_6')
// (11, 13, 'sp4_r_v_b_7')
// (12, 9, 'sp12_h_r_6')
// (12, 9, 'sp4_h_l_39')
// (12, 9, 'sp4_h_r_15')
// (12, 9, 'sp4_v_t_42')
// (12, 10, 'local_g2_2')
// (12, 10, 'lutff_1/in_3')
// (12, 10, 'lutff_7/in_3')
// (12, 10, 'sp4_v_b_42')
// (12, 11, 'sp4_v_b_31')
// (12, 12, 'sp4_h_r_19')
// (12, 12, 'sp4_v_b_18')
// (12, 13, 'sp4_v_b_7')
// (13, 9, 'sp12_h_r_9')
// (13, 9, 'sp4_h_r_26')
// (13, 12, 'sp4_h_r_30')
// (14, 9, 'local_g0_2')
// (14, 9, 'lutff_0/in_0')
// (14, 9, 'lutff_3/in_3')
// (14, 9, 'sp12_h_r_10')
// (14, 9, 'sp4_h_r_39')
// (14, 10, 'sp4_r_v_b_39')
// (14, 11, 'sp4_r_v_b_26')
// (14, 12, 'local_g2_3')
// (14, 12, 'local_g3_3')
// (14, 12, 'lutff_0/in_1')
// (14, 12, 'lutff_2/in_0')
// (14, 12, 'sp4_h_r_43')
// (14, 12, 'sp4_r_v_b_15')
// (14, 13, 'sp4_r_v_b_2')
// (15, 9, 'sp12_h_r_13')
// (15, 9, 'sp4_h_l_39')
// (15, 9, 'sp4_v_t_39')
// (15, 10, 'sp4_v_b_39')
// (15, 11, 'sp4_v_b_26')
// (15, 12, 'local_g0_7')
// (15, 12, 'local_g1_7')
// (15, 12, 'lutff_2/in_0')
// (15, 12, 'lutff_4/in_1')
// (15, 12, 'sp4_h_l_43')
// (15, 12, 'sp4_v_b_15')
// (15, 13, 'sp4_v_b_2')
// (16, 9, 'sp12_h_r_14')
// (17, 9, 'sp12_h_r_17')
// (18, 9, 'sp12_h_r_18')
// (19, 9, 'sp12_h_r_21')
// (20, 9, 'sp12_h_r_22')
// (21, 9, 'sp12_h_l_22')

wire n153;
// (8, 10, 'neigh_op_tnr_3')
// (8, 11, 'neigh_op_rgt_3')
// (8, 12, 'neigh_op_bnr_3')
// (9, 10, 'neigh_op_top_3')
// (9, 11, 'lutff_3/out')
// (9, 11, 'sp4_r_v_b_39')
// (9, 12, 'neigh_op_bot_3')
// (9, 12, 'sp4_r_v_b_26')
// (9, 13, 'sp4_r_v_b_15')
// (9, 14, 'sp4_r_v_b_2')
// (9, 15, 'sp4_r_v_b_39')
// (9, 16, 'sp4_r_v_b_26')
// (9, 17, 'sp4_r_v_b_15')
// (9, 18, 'sp4_r_v_b_2')
// (10, 10, 'neigh_op_tnl_3')
// (10, 10, 'sp4_v_t_39')
// (10, 11, 'neigh_op_lft_3')
// (10, 11, 'sp4_v_b_39')
// (10, 12, 'neigh_op_bnl_3')
// (10, 12, 'sp4_v_b_26')
// (10, 13, 'sp4_v_b_15')
// (10, 14, 'sp4_v_b_2')
// (10, 14, 'sp4_v_t_39')
// (10, 15, 'sp4_v_b_39')
// (10, 16, 'sp4_v_b_26')
// (10, 17, 'sp4_v_b_15')
// (10, 18, 'local_g0_2')
// (10, 18, 'lutff_global/cen')
// (10, 18, 'sp4_v_b_2')

reg n154 = 0;
// (8, 11, 'neigh_op_tnr_1')
// (8, 11, 'sp4_r_v_b_47')
// (8, 12, 'neigh_op_rgt_1')
// (8, 12, 'sp4_r_v_b_34')
// (8, 13, 'neigh_op_bnr_1')
// (8, 13, 'sp4_r_v_b_23')
// (8, 14, 'sp4_r_v_b_10')
// (9, 10, 'sp4_h_r_10')
// (9, 10, 'sp4_v_t_47')
// (9, 11, 'neigh_op_top_1')
// (9, 11, 'sp4_v_b_47')
// (9, 12, 'local_g0_1')
// (9, 12, 'lutff_1/in_0')
// (9, 12, 'lutff_1/out')
// (9, 12, 'sp4_v_b_34')
// (9, 13, 'neigh_op_bot_1')
// (9, 13, 'sp4_v_b_23')
// (9, 14, 'sp4_v_b_10')
// (10, 10, 'sp4_h_r_23')
// (10, 11, 'neigh_op_tnl_1')
// (10, 12, 'neigh_op_lft_1')
// (10, 13, 'neigh_op_bnl_1')
// (11, 10, 'local_g2_2')
// (11, 10, 'local_g3_2')
// (11, 10, 'lutff_0/in_1')
// (11, 10, 'lutff_1/in_1')
// (11, 10, 'lutff_7/in_1')
// (11, 10, 'sp4_h_r_34')
// (12, 10, 'sp4_h_r_47')
// (13, 10, 'sp4_h_l_47')

wire n155;
// (8, 11, 'neigh_op_tnr_4')
// (8, 12, 'neigh_op_rgt_4')
// (8, 13, 'neigh_op_bnr_4')
// (9, 11, 'neigh_op_top_4')
// (9, 12, 'local_g0_4')
// (9, 12, 'lutff_1/in_3')
// (9, 12, 'lutff_3/in_3')
// (9, 12, 'lutff_4/out')
// (9, 12, 'lutff_7/in_3')
// (9, 13, 'neigh_op_bot_4')
// (10, 11, 'neigh_op_tnl_4')
// (10, 12, 'neigh_op_lft_4')
// (10, 13, 'neigh_op_bnl_4')

wire n156;
// (8, 11, 'neigh_op_tnr_5')
// (8, 12, 'neigh_op_rgt_5')
// (8, 12, 'sp4_r_v_b_42')
// (8, 13, 'neigh_op_bnr_5')
// (8, 13, 'sp4_r_v_b_31')
// (8, 14, 'sp4_r_v_b_18')
// (8, 15, 'sp4_r_v_b_7')
// (9, 11, 'neigh_op_top_5')
// (9, 11, 'sp4_v_t_42')
// (9, 12, 'lutff_5/out')
// (9, 12, 'sp4_v_b_42')
// (9, 13, 'neigh_op_bot_5')
// (9, 13, 'sp4_v_b_31')
// (9, 14, 'local_g0_2')
// (9, 14, 'lutff_7/in_3')
// (9, 14, 'sp4_v_b_18')
// (9, 15, 'sp4_v_b_7')
// (10, 11, 'neigh_op_tnl_5')
// (10, 12, 'neigh_op_lft_5')
// (10, 13, 'neigh_op_bnl_5')

wire n157;
// (8, 12, 'sp12_h_r_1')
// (9, 12, 'sp12_h_r_2')
// (10, 12, 'sp12_h_r_5')
// (11, 12, 'sp12_h_r_6')
// (12, 12, 'sp12_h_r_9')
// (13, 12, 'sp12_h_r_10')
// (14, 12, 'local_g1_5')
// (14, 12, 'lutff_5/in_3')
// (14, 12, 'sp12_h_r_13')
// (15, 12, 'sp12_h_r_14')
// (15, 20, 'sp4_h_r_6')
// (16, 12, 'sp12_h_r_17')
// (16, 20, 'local_g1_3')
// (16, 20, 'lutff_1/in_1')
// (16, 20, 'sp4_h_r_19')
// (17, 12, 'sp12_h_r_18')
// (17, 20, 'sp4_h_r_30')
// (18, 11, 'neigh_op_tnr_7')
// (18, 12, 'neigh_op_rgt_7')
// (18, 12, 'sp12_h_r_21')
// (18, 13, 'neigh_op_bnr_7')
// (18, 17, 'sp4_r_v_b_36')
// (18, 18, 'sp4_r_v_b_25')
// (18, 19, 'sp4_r_v_b_12')
// (18, 20, 'sp4_h_r_43')
// (18, 20, 'sp4_r_v_b_1')
// (19, 7, 'sp12_v_t_22')
// (19, 8, 'sp12_v_b_22')
// (19, 9, 'sp12_v_b_21')
// (19, 10, 'sp12_v_b_18')
// (19, 11, 'neigh_op_top_7')
// (19, 11, 'sp12_v_b_17')
// (19, 12, 'lutff_7/out')
// (19, 12, 'sp12_h_r_22')
// (19, 12, 'sp12_v_b_14')
// (19, 13, 'neigh_op_bot_7')
// (19, 13, 'sp12_v_b_13')
// (19, 14, 'sp12_v_b_10')
// (19, 15, 'sp12_v_b_9')
// (19, 16, 'sp12_v_b_6')
// (19, 16, 'sp4_v_t_36')
// (19, 17, 'sp12_v_b_5')
// (19, 17, 'sp4_v_b_36')
// (19, 18, 'sp12_v_b_2')
// (19, 18, 'sp4_v_b_25')
// (19, 19, 'sp12_v_b_1')
// (19, 19, 'sp4_v_b_12')
// (19, 20, 'local_g0_1')
// (19, 20, 'lutff_6/in_1')
// (19, 20, 'sp4_h_l_43')
// (19, 20, 'sp4_v_b_1')
// (20, 11, 'neigh_op_tnl_7')
// (20, 12, 'neigh_op_lft_7')
// (20, 12, 'sp12_h_l_22')
// (20, 13, 'neigh_op_bnl_7')

reg n158 = 0;
// (8, 13, 'sp4_r_v_b_39')
// (8, 14, 'sp4_r_v_b_26')
// (8, 15, 'sp4_r_v_b_15')
// (8, 16, 'sp4_r_v_b_2')
// (9, 12, 'sp4_h_r_2')
// (9, 12, 'sp4_v_t_39')
// (9, 13, 'sp4_v_b_39')
// (9, 14, 'sp4_v_b_26')
// (9, 15, 'sp4_v_b_15')
// (9, 16, 'local_g1_2')
// (9, 16, 'lutff_7/in_0')
// (9, 16, 'sp4_r_v_b_42')
// (9, 16, 'sp4_v_b_2')
// (9, 17, 'sp4_r_v_b_31')
// (9, 18, 'local_g3_2')
// (9, 18, 'lutff_1/in_0')
// (9, 18, 'sp4_r_v_b_18')
// (9, 19, 'sp4_r_v_b_7')
// (10, 11, 'neigh_op_tnr_5')
// (10, 12, 'neigh_op_rgt_5')
// (10, 12, 'sp12_h_r_1')
// (10, 12, 'sp12_v_t_22')
// (10, 12, 'sp4_h_r_15')
// (10, 13, 'neigh_op_bnr_5')
// (10, 13, 'sp12_v_b_22')
// (10, 14, 'sp12_v_b_21')
// (10, 15, 'sp12_v_b_18')
// (10, 15, 'sp4_v_t_42')
// (10, 16, 'sp12_v_b_17')
// (10, 16, 'sp4_v_b_42')
// (10, 17, 'sp12_v_b_14')
// (10, 17, 'sp4_v_b_31')
// (10, 18, 'sp12_v_b_13')
// (10, 18, 'sp4_v_b_18')
// (10, 19, 'local_g2_2')
// (10, 19, 'lutff_5/in_3')
// (10, 19, 'sp12_v_b_10')
// (10, 19, 'sp4_h_r_7')
// (10, 19, 'sp4_v_b_7')
// (10, 20, 'local_g3_1')
// (10, 20, 'lutff_3/in_3')
// (10, 20, 'sp12_v_b_9')
// (10, 21, 'sp12_v_b_6')
// (10, 22, 'sp12_v_b_5')
// (10, 23, 'sp12_v_b_2')
// (10, 24, 'sp12_h_r_1')
// (10, 24, 'sp12_v_b_1')
// (11, 5, 'sp12_v_t_22')
// (11, 6, 'sp12_v_b_22')
// (11, 7, 'sp12_v_b_21')
// (11, 8, 'sp12_v_b_18')
// (11, 9, 'sp12_v_b_17')
// (11, 10, 'sp12_v_b_14')
// (11, 11, 'neigh_op_top_5')
// (11, 11, 'sp12_v_b_13')
// (11, 12, 'lutff_5/out')
// (11, 12, 'sp12_h_r_2')
// (11, 12, 'sp12_v_b_10')
// (11, 12, 'sp4_h_r_26')
// (11, 13, 'local_g1_5')
// (11, 13, 'lutff_3/in_3')
// (11, 13, 'neigh_op_bot_5')
// (11, 13, 'sp12_v_b_9')
// (11, 14, 'sp12_v_b_6')
// (11, 15, 'sp12_v_b_5')
// (11, 16, 'sp12_v_b_2')
// (11, 17, 'sp12_v_b_1')
// (11, 17, 'sp12_v_t_22')
// (11, 18, 'sp12_v_b_22')
// (11, 19, 'sp12_v_b_21')
// (11, 19, 'sp4_h_r_18')
// (11, 20, 'sp12_v_b_18')
// (11, 21, 'sp12_v_b_17')
// (11, 22, 'local_g3_6')
// (11, 22, 'lutff_5/in_0')
// (11, 22, 'sp12_v_b_14')
// (11, 23, 'sp12_v_b_13')
// (11, 24, 'sp12_h_r_2')
// (11, 24, 'sp12_v_b_10')
// (11, 25, 'sp12_v_b_9')
// (11, 26, 'sp12_v_b_6')
// (11, 27, 'sp12_v_b_5')
// (11, 28, 'sp12_v_b_2')
// (11, 29, 'sp12_v_b_1')
// (12, 11, 'neigh_op_tnl_5')
// (12, 12, 'neigh_op_lft_5')
// (12, 12, 'sp12_h_r_5')
// (12, 12, 'sp4_h_r_39')
// (12, 13, 'local_g3_5')
// (12, 13, 'lutff_5/in_3')
// (12, 13, 'neigh_op_bnl_5')
// (12, 19, 'local_g3_7')
// (12, 19, 'lutff_5/in_3')
// (12, 19, 'sp4_h_r_31')
// (12, 20, 'local_g1_1')
// (12, 20, 'lutff_5/in_3')
// (12, 20, 'sp4_h_r_1')
// (12, 24, 'sp12_h_r_5')
// (13, 12, 'sp12_h_r_6')
// (13, 12, 'sp4_h_l_39')
// (13, 13, 'sp4_r_v_b_41')
// (13, 14, 'sp4_r_v_b_28')
// (13, 15, 'sp4_r_v_b_17')
// (13, 16, 'local_g1_4')
// (13, 16, 'lutff_3/in_0')
// (13, 16, 'sp4_r_v_b_4')
// (13, 19, 'sp4_h_r_42')
// (13, 20, 'sp4_h_r_12')
// (13, 20, 'sp4_r_v_b_37')
// (13, 21, 'sp4_r_v_b_24')
// (13, 22, 'sp4_r_v_b_13')
// (13, 23, 'sp4_r_v_b_0')
// (13, 24, 'sp12_h_r_6')
// (14, 12, 'sp12_h_r_9')
// (14, 12, 'sp4_h_r_4')
// (14, 12, 'sp4_v_t_41')
// (14, 13, 'local_g3_1')
// (14, 13, 'lutff_5/in_3')
// (14, 13, 'sp4_v_b_41')
// (14, 14, 'sp4_v_b_28')
// (14, 15, 'sp4_v_b_17')
// (14, 16, 'sp4_v_b_4')
// (14, 19, 'sp4_h_l_42')
// (14, 19, 'sp4_h_r_10')
// (14, 19, 'sp4_v_t_37')
// (14, 20, 'sp4_h_r_25')
// (14, 20, 'sp4_v_b_37')
// (14, 21, 'sp4_h_r_4')
// (14, 21, 'sp4_v_b_24')
// (14, 22, 'local_g1_5')
// (14, 22, 'lutff_3/in_3')
// (14, 22, 'sp4_v_b_13')
// (14, 23, 'sp4_v_b_0')
// (14, 24, 'sp12_h_r_9')
// (15, 9, 'sp4_r_v_b_45')
// (15, 10, 'sp4_r_v_b_32')
// (15, 11, 'sp4_r_v_b_21')
// (15, 12, 'sp12_h_r_10')
// (15, 12, 'sp4_h_r_17')
// (15, 12, 'sp4_r_v_b_8')
// (15, 13, 'sp4_r_v_b_37')
// (15, 14, 'sp4_r_v_b_24')
// (15, 15, 'local_g2_5')
// (15, 15, 'lutff_5/in_0')
// (15, 15, 'sp4_r_v_b_13')
// (15, 16, 'sp4_r_v_b_0')
// (15, 17, 'local_g3_5')
// (15, 17, 'lutff_5/in_3')
// (15, 17, 'sp4_r_v_b_45')
// (15, 18, 'local_g2_0')
// (15, 18, 'lutff_5/in_3')
// (15, 18, 'sp4_r_v_b_32')
// (15, 19, 'local_g3_5')
// (15, 19, 'lutff_5/in_3')
// (15, 19, 'sp4_h_r_23')
// (15, 19, 'sp4_r_v_b_21')
// (15, 20, 'sp4_h_r_36')
// (15, 20, 'sp4_r_v_b_8')
// (15, 21, 'sp4_h_r_17')
// (15, 24, 'sp12_h_r_10')
// (16, 8, 'sp4_v_t_45')
// (16, 9, 'sp4_v_b_45')
// (16, 10, 'sp4_v_b_32')
// (16, 11, 'local_g1_5')
// (16, 11, 'lutff_5/in_3')
// (16, 11, 'sp4_v_b_21')
// (16, 12, 'sp12_h_r_13')
// (16, 12, 'sp4_h_r_28')
// (16, 12, 'sp4_h_r_6')
// (16, 12, 'sp4_v_b_8')
// (16, 12, 'sp4_v_t_37')
// (16, 13, 'sp4_v_b_37')
// (16, 14, 'local_g2_0')
// (16, 14, 'lutff_3/in_1')
// (16, 14, 'sp4_v_b_24')
// (16, 15, 'sp4_v_b_13')
// (16, 16, 'local_g0_0')
// (16, 16, 'lutff_5/in_1')
// (16, 16, 'sp4_v_b_0')
// (16, 16, 'sp4_v_t_45')
// (16, 17, 'local_g3_5')
// (16, 17, 'lutff_5/in_3')
// (16, 17, 'sp4_v_b_45')
// (16, 18, 'local_g2_0')
// (16, 18, 'lutff_5/in_3')
// (16, 18, 'sp4_v_b_32')
// (16, 19, 'local_g1_5')
// (16, 19, 'lutff_3/in_3')
// (16, 19, 'sp4_h_r_34')
// (16, 19, 'sp4_v_b_21')
// (16, 20, 'sp4_h_l_36')
// (16, 20, 'sp4_v_b_8')
// (16, 21, 'local_g2_4')
// (16, 21, 'lutff_3/in_3')
// (16, 21, 'sp4_h_r_28')
// (16, 24, 'sp12_h_r_13')
// (17, 9, 'sp4_r_v_b_47')
// (17, 10, 'sp4_r_v_b_34')
// (17, 11, 'local_g3_7')
// (17, 11, 'lutff_6/in_0')
// (17, 11, 'sp4_r_v_b_23')
// (17, 12, 'sp12_h_r_14')
// (17, 12, 'sp4_h_r_19')
// (17, 12, 'sp4_h_r_41')
// (17, 12, 'sp4_r_v_b_10')
// (17, 13, 'sp4_r_v_b_47')
// (17, 14, 'local_g2_2')
// (17, 14, 'lutff_2/in_0')
// (17, 14, 'sp4_r_v_b_34')
// (17, 15, 'sp4_r_v_b_23')
// (17, 16, 'sp4_r_v_b_10')
// (17, 16, 'sp4_r_v_b_41')
// (17, 17, 'sp4_r_v_b_28')
// (17, 18, 'sp4_r_v_b_17')
// (17, 19, 'sp4_h_r_47')
// (17, 19, 'sp4_r_v_b_4')
// (17, 21, 'sp4_h_r_41')
// (17, 24, 'sp12_h_r_14')
// (18, 8, 'sp4_v_t_47')
// (18, 9, 'sp4_v_b_47')
// (18, 10, 'sp4_v_b_34')
// (18, 11, 'sp4_v_b_23')
// (18, 12, 'local_g1_1')
// (18, 12, 'lutff_5/in_3')
// (18, 12, 'sp12_h_r_17')
// (18, 12, 'sp4_h_l_41')
// (18, 12, 'sp4_h_r_30')
// (18, 12, 'sp4_h_r_4')
// (18, 12, 'sp4_v_b_10')
// (18, 12, 'sp4_v_t_47')
// (18, 13, 'sp4_v_b_47')
// (18, 14, 'sp4_v_b_34')
// (18, 15, 'sp4_v_b_23')
// (18, 15, 'sp4_v_t_41')
// (18, 16, 'sp4_v_b_10')
// (18, 16, 'sp4_v_b_41')
// (18, 17, 'sp4_v_b_28')
// (18, 18, 'local_g1_1')
// (18, 18, 'lutff_3/in_3')
// (18, 18, 'sp4_v_b_17')
// (18, 19, 'sp4_h_l_47')
// (18, 19, 'sp4_h_r_1')
// (18, 19, 'sp4_v_b_4')
// (18, 21, 'sp4_h_l_41')
// (18, 21, 'sp4_h_r_1')
// (18, 24, 'sp12_h_r_17')
// (19, 9, 'sp4_r_v_b_37')
// (19, 10, 'local_g0_0')
// (19, 10, 'lutff_5/in_1')
// (19, 10, 'sp4_r_v_b_24')
// (19, 11, 'local_g2_5')
// (19, 11, 'lutff_5/in_0')
// (19, 11, 'sp4_r_v_b_13')
// (19, 12, 'sp12_h_r_18')
// (19, 12, 'sp4_h_r_17')
// (19, 12, 'sp4_h_r_43')
// (19, 12, 'sp4_r_v_b_0')
// (19, 13, 'sp4_r_v_b_43')
// (19, 14, 'local_g0_6')
// (19, 14, 'lutff_0/in_0')
// (19, 14, 'sp4_r_v_b_30')
// (19, 15, 'sp4_r_v_b_19')
// (19, 16, 'local_g1_6')
// (19, 16, 'lutff_5/in_0')
// (19, 16, 'sp4_r_v_b_6')
// (19, 17, 'sp4_r_v_b_39')
// (19, 18, 'sp4_r_v_b_26')
// (19, 19, 'local_g1_4')
// (19, 19, 'lutff_4/in_3')
// (19, 19, 'sp4_h_r_12')
// (19, 19, 'sp4_r_v_b_15')
// (19, 20, 'sp4_r_v_b_2')
// (19, 21, 'sp4_h_r_12')
// (19, 24, 'sp12_h_r_18')
// (19, 25, 'sp4_r_v_b_41')
// (19, 26, 'sp4_r_v_b_28')
// (19, 27, 'sp4_r_v_b_17')
// (19, 28, 'sp4_r_v_b_4')
// (20, 8, 'sp4_v_t_37')
// (20, 9, 'sp4_v_b_37')
// (20, 10, 'sp4_v_b_24')
// (20, 11, 'local_g0_5')
// (20, 11, 'lutff_4/in_3')
// (20, 11, 'sp4_v_b_13')
// (20, 12, 'local_g1_5')
// (20, 12, 'lutff_5/in_3')
// (20, 12, 'sp12_h_r_21')
// (20, 12, 'sp4_h_l_43')
// (20, 12, 'sp4_h_r_28')
// (20, 12, 'sp4_h_r_9')
// (20, 12, 'sp4_v_b_0')
// (20, 12, 'sp4_v_t_43')
// (20, 13, 'sp4_v_b_43')
// (20, 14, 'sp4_v_b_30')
// (20, 15, 'sp4_v_b_19')
// (20, 16, 'local_g0_6')
// (20, 16, 'lutff_5/in_3')
// (20, 16, 'sp4_v_b_6')
// (20, 16, 'sp4_v_t_39')
// (20, 17, 'sp4_v_b_39')
// (20, 18, 'sp4_v_b_26')
// (20, 19, 'local_g1_7')
// (20, 19, 'lutff_5/in_3')
// (20, 19, 'sp4_h_r_25')
// (20, 19, 'sp4_v_b_15')
// (20, 20, 'local_g0_2')
// (20, 20, 'lutff_5/in_3')
// (20, 20, 'sp4_v_b_2')
// (20, 21, 'local_g3_1')
// (20, 21, 'lutff_5/in_3')
// (20, 21, 'sp4_h_r_25')
// (20, 24, 'sp12_h_r_21')
// (20, 24, 'sp4_h_r_10')
// (20, 24, 'sp4_v_t_41')
// (20, 25, 'sp4_v_b_41')
// (20, 26, 'local_g3_4')
// (20, 26, 'lutff_2/in_3')
// (20, 26, 'sp4_v_b_28')
// (20, 27, 'sp4_v_b_17')
// (20, 28, 'sp4_v_b_4')
// (21, 9, 'sp4_r_v_b_41')
// (21, 10, 'sp4_r_v_b_28')
// (21, 11, 'local_g3_1')
// (21, 11, 'lutff_5/in_3')
// (21, 11, 'sp4_r_v_b_17')
// (21, 12, 'local_g0_6')
// (21, 12, 'lutff_5/in_3')
// (21, 12, 'sp12_h_r_22')
// (21, 12, 'sp4_h_r_20')
// (21, 12, 'sp4_h_r_41')
// (21, 12, 'sp4_r_v_b_4')
// (21, 16, 'sp4_r_v_b_41')
// (21, 17, 'local_g0_4')
// (21, 17, 'lutff_5/in_3')
// (21, 17, 'sp4_r_v_b_28')
// (21, 18, 'sp4_r_v_b_17')
// (21, 19, 'sp4_h_r_36')
// (21, 19, 'sp4_r_v_b_4')
// (21, 20, 'local_g2_6')
// (21, 20, 'lutff_5/in_3')
// (21, 20, 'sp4_r_v_b_38')
// (21, 21, 'sp4_h_r_36')
// (21, 21, 'sp4_r_v_b_27')
// (21, 22, 'sp4_r_v_b_14')
// (21, 22, 'sp4_r_v_b_36')
// (21, 23, 'sp4_r_v_b_25')
// (21, 23, 'sp4_r_v_b_3')
// (21, 24, 'local_g0_6')
// (21, 24, 'lutff_1/in_3')
// (21, 24, 'sp12_h_r_22')
// (21, 24, 'sp4_h_r_23')
// (21, 24, 'sp4_r_v_b_12')
// (21, 25, 'sp4_r_v_b_1')
// (22, 8, 'sp4_v_t_41')
// (22, 9, 'sp4_v_b_41')
// (22, 10, 'sp4_v_b_28')
// (22, 11, 'sp4_v_b_17')
// (22, 12, 'local_g3_1')
// (22, 12, 'lutff_5/in_3')
// (22, 12, 'sp12_h_l_22')
// (22, 12, 'sp12_v_t_22')
// (22, 12, 'sp4_h_l_41')
// (22, 12, 'sp4_h_r_33')
// (22, 12, 'sp4_v_b_4')
// (22, 13, 'sp12_v_b_22')
// (22, 14, 'local_g3_5')
// (22, 14, 'lutff_5/in_3')
// (22, 14, 'sp12_v_b_21')
// (22, 15, 'sp12_v_b_18')
// (22, 15, 'sp4_v_t_41')
// (22, 16, 'sp12_v_b_17')
// (22, 16, 'sp4_v_b_41')
// (22, 17, 'sp12_v_b_14')
// (22, 17, 'sp4_v_b_28')
// (22, 18, 'sp12_v_b_13')
// (22, 18, 'sp4_v_b_17')
// (22, 19, 'local_g2_2')
// (22, 19, 'lutff_3/in_3')
// (22, 19, 'sp12_v_b_10')
// (22, 19, 'sp4_h_l_36')
// (22, 19, 'sp4_h_r_4')
// (22, 19, 'sp4_v_b_4')
// (22, 19, 'sp4_v_t_38')
// (22, 20, 'sp12_v_b_9')
// (22, 20, 'sp4_v_b_38')
// (22, 21, 'local_g3_6')
// (22, 21, 'lutff_5/in_0')
// (22, 21, 'sp12_v_b_6')
// (22, 21, 'sp4_h_l_36')
// (22, 21, 'sp4_v_b_27')
// (22, 21, 'sp4_v_t_36')
// (22, 22, 'sp12_v_b_5')
// (22, 22, 'sp4_v_b_14')
// (22, 22, 'sp4_v_b_36')
// (22, 23, 'local_g2_2')
// (22, 23, 'lutff_5/in_3')
// (22, 23, 'sp12_v_b_2')
// (22, 23, 'sp4_v_b_25')
// (22, 23, 'sp4_v_b_3')
// (22, 24, 'sp12_h_l_22')
// (22, 24, 'sp12_v_b_1')
// (22, 24, 'sp4_h_r_34')
// (22, 24, 'sp4_v_b_12')
// (22, 25, 'sp4_v_b_1')
// (23, 12, 'local_g2_4')
// (23, 12, 'lutff_5/in_3')
// (23, 12, 'sp4_h_r_44')
// (23, 13, 'local_g3_4')
// (23, 13, 'lutff_3/in_0')
// (23, 13, 'sp4_r_v_b_44')
// (23, 14, 'local_g0_2')
// (23, 14, 'lutff_5/in_3')
// (23, 14, 'sp4_r_v_b_33')
// (23, 15, 'local_g3_4')
// (23, 15, 'lutff_5/in_0')
// (23, 15, 'sp4_r_v_b_20')
// (23, 16, 'local_g2_1')
// (23, 16, 'lutff_5/in_0')
// (23, 16, 'sp4_r_v_b_9')
// (23, 17, 'sp4_r_v_b_37')
// (23, 18, 'sp4_r_v_b_24')
// (23, 19, 'sp4_h_r_17')
// (23, 19, 'sp4_r_v_b_13')
// (23, 20, 'local_g1_0')
// (23, 20, 'lutff_5/in_0')
// (23, 20, 'sp4_r_v_b_0')
// (23, 24, 'sp4_h_r_47')
// (24, 12, 'sp4_h_l_44')
// (24, 12, 'sp4_v_t_44')
// (24, 13, 'local_g2_4')
// (24, 13, 'lutff_1/in_3')
// (24, 13, 'sp4_v_b_44')
// (24, 14, 'local_g2_1')
// (24, 14, 'lutff_5/in_0')
// (24, 14, 'sp4_v_b_33')
// (24, 15, 'sp4_v_b_20')
// (24, 16, 'local_g1_1')
// (24, 16, 'lutff_1/in_3')
// (24, 16, 'sp4_v_b_9')
// (24, 16, 'sp4_v_t_37')
// (24, 17, 'local_g3_5')
// (24, 17, 'lutff_5/in_3')
// (24, 17, 'sp4_v_b_37')
// (24, 18, 'sp4_v_b_24')
// (24, 19, 'sp4_h_r_28')
// (24, 19, 'sp4_v_b_13')
// (24, 20, 'sp4_v_b_0')
// (24, 24, 'sp4_h_l_47')
// (25, 19, 'sp4_h_r_41')
// (26, 19, 'sp4_h_l_41')

reg n159 = 0;
// (8, 13, 'sp4_r_v_b_45')
// (8, 14, 'sp4_r_v_b_32')
// (8, 15, 'sp4_r_v_b_21')
// (8, 16, 'sp4_r_v_b_8')
// (8, 17, 'sp4_r_v_b_45')
// (8, 18, 'sp4_r_v_b_32')
// (8, 19, 'sp4_r_v_b_21')
// (8, 20, 'sp4_r_v_b_8')
// (9, 12, 'sp4_h_r_8')
// (9, 12, 'sp4_v_t_45')
// (9, 13, 'sp4_v_b_45')
// (9, 14, 'sp4_v_b_32')
// (9, 15, 'local_g1_5')
// (9, 15, 'lutff_5/in_3')
// (9, 15, 'sp4_v_b_21')
// (9, 16, 'sp4_v_b_8')
// (9, 16, 'sp4_v_t_45')
// (9, 17, 'local_g3_5')
// (9, 17, 'lutff_1/in_3')
// (9, 17, 'sp4_v_b_45')
// (9, 18, 'sp4_v_b_32')
// (9, 19, 'sp4_v_b_21')
// (9, 20, 'sp4_v_b_8')
// (10, 11, 'neigh_op_tnr_0')
// (10, 12, 'neigh_op_rgt_0')
// (10, 12, 'sp4_h_r_21')
// (10, 12, 'sp4_h_r_5')
// (10, 13, 'neigh_op_bnr_0')
// (10, 17, 'sp4_r_v_b_37')
// (10, 18, 'sp4_r_v_b_24')
// (10, 19, 'local_g2_5')
// (10, 19, 'lutff_0/in_3')
// (10, 19, 'sp4_r_v_b_13')
// (10, 20, 'local_g1_0')
// (10, 20, 'lutff_6/in_3')
// (10, 20, 'sp4_r_v_b_0')
// (11, 8, 'sp12_v_t_23')
// (11, 9, 'sp12_v_b_23')
// (11, 10, 'sp12_v_b_20')
// (11, 10, 'sp4_r_v_b_41')
// (11, 11, 'neigh_op_top_0')
// (11, 11, 'sp12_v_b_19')
// (11, 11, 'sp4_r_v_b_28')
// (11, 11, 'sp4_r_v_b_44')
// (11, 12, 'lutff_0/out')
// (11, 12, 'sp12_v_b_16')
// (11, 12, 'sp4_h_r_16')
// (11, 12, 'sp4_h_r_32')
// (11, 12, 'sp4_r_v_b_17')
// (11, 12, 'sp4_r_v_b_33')
// (11, 13, 'local_g1_0')
// (11, 13, 'lutff_6/in_3')
// (11, 13, 'neigh_op_bot_0')
// (11, 13, 'sp12_v_b_15')
// (11, 13, 'sp4_r_v_b_20')
// (11, 13, 'sp4_r_v_b_4')
// (11, 14, 'sp12_v_b_12')
// (11, 14, 'sp4_r_v_b_9')
// (11, 15, 'sp12_v_b_11')
// (11, 16, 'sp12_v_b_8')
// (11, 16, 'sp4_v_t_37')
// (11, 17, 'sp12_v_b_7')
// (11, 17, 'sp4_v_b_37')
// (11, 18, 'sp12_v_b_4')
// (11, 18, 'sp4_v_b_24')
// (11, 19, 'sp12_v_b_3')
// (11, 19, 'sp4_v_b_13')
// (11, 20, 'sp12_h_r_0')
// (11, 20, 'sp12_v_b_0')
// (11, 20, 'sp12_v_t_23')
// (11, 20, 'sp4_v_b_0')
// (11, 21, 'sp12_v_b_23')
// (11, 22, 'local_g3_4')
// (11, 22, 'lutff_0/in_3')
// (11, 22, 'sp12_v_b_20')
// (11, 23, 'sp12_v_b_19')
// (11, 24, 'sp12_v_b_16')
// (11, 25, 'sp12_v_b_15')
// (11, 26, 'sp12_v_b_12')
// (11, 27, 'sp12_v_b_11')
// (11, 28, 'sp12_v_b_8')
// (11, 29, 'sp12_v_b_7')
// (11, 30, 'sp12_v_b_4')
// (11, 31, 'sp12_v_b_3')
// (11, 32, 'sp12_v_b_0')
// (12, 9, 'sp4_v_t_41')
// (12, 10, 'sp4_v_b_41')
// (12, 10, 'sp4_v_t_44')
// (12, 11, 'neigh_op_tnl_0')
// (12, 11, 'sp4_v_b_28')
// (12, 11, 'sp4_v_b_44')
// (12, 12, 'neigh_op_lft_0')
// (12, 12, 'sp4_h_r_29')
// (12, 12, 'sp4_h_r_45')
// (12, 12, 'sp4_v_b_17')
// (12, 12, 'sp4_v_b_33')
// (12, 13, 'local_g3_0')
// (12, 13, 'lutff_0/in_3')
// (12, 13, 'neigh_op_bnl_0')
// (12, 13, 'sp4_h_r_10')
// (12, 13, 'sp4_r_v_b_36')
// (12, 13, 'sp4_v_b_20')
// (12, 13, 'sp4_v_b_4')
// (12, 14, 'sp4_h_r_9')
// (12, 14, 'sp4_r_v_b_25')
// (12, 14, 'sp4_v_b_9')
// (12, 15, 'sp4_r_v_b_12')
// (12, 16, 'sp4_r_v_b_1')
// (12, 17, 'sp4_r_v_b_44')
// (12, 18, 'sp4_r_v_b_33')
// (12, 19, 'local_g3_4')
// (12, 19, 'lutff_0/in_3')
// (12, 19, 'sp4_r_v_b_20')
// (12, 20, 'local_g2_1')
// (12, 20, 'lutff_0/in_3')
// (12, 20, 'sp12_h_r_3')
// (12, 20, 'sp4_r_v_b_9')
// (13, 12, 'sp4_h_l_45')
// (13, 12, 'sp4_h_r_11')
// (13, 12, 'sp4_h_r_4')
// (13, 12, 'sp4_h_r_40')
// (13, 12, 'sp4_v_t_36')
// (13, 13, 'sp4_h_r_23')
// (13, 13, 'sp4_v_b_36')
// (13, 14, 'sp4_h_r_20')
// (13, 14, 'sp4_v_b_25')
// (13, 15, 'sp4_v_b_12')
// (13, 16, 'local_g0_1')
// (13, 16, 'lutff_6/in_1')
// (13, 16, 'sp4_v_b_1')
// (13, 16, 'sp4_v_t_44')
// (13, 17, 'sp4_v_b_44')
// (13, 18, 'sp4_v_b_33')
// (13, 19, 'sp4_v_b_20')
// (13, 20, 'sp12_h_r_4')
// (13, 20, 'sp4_v_b_9')
// (13, 21, 'sp4_r_v_b_40')
// (13, 22, 'sp4_r_v_b_29')
// (13, 23, 'sp4_r_v_b_16')
// (13, 24, 'sp4_r_v_b_5')
// (14, 12, 'local_g1_6')
// (14, 12, 'lutff_6/in_1')
// (14, 12, 'sp4_h_l_40')
// (14, 12, 'sp4_h_r_1')
// (14, 12, 'sp4_h_r_17')
// (14, 12, 'sp4_h_r_22')
// (14, 12, 'sp4_h_r_5')
// (14, 13, 'local_g3_2')
// (14, 13, 'lutff_0/in_3')
// (14, 13, 'sp4_h_r_34')
// (14, 14, 'sp4_h_r_33')
// (14, 20, 'sp12_h_r_7')
// (14, 20, 'sp4_h_r_5')
// (14, 20, 'sp4_v_t_40')
// (14, 21, 'sp4_v_b_40')
// (14, 22, 'local_g2_5')
// (14, 22, 'lutff_0/in_3')
// (14, 22, 'sp4_v_b_29')
// (14, 23, 'sp4_v_b_16')
// (14, 24, 'sp4_v_b_5')
// (15, 10, 'sp4_r_v_b_41')
// (15, 11, 'sp4_r_v_b_28')
// (15, 12, 'local_g2_3')
// (15, 12, 'lutff_0/in_1')
// (15, 12, 'sp4_h_r_12')
// (15, 12, 'sp4_h_r_16')
// (15, 12, 'sp4_h_r_28')
// (15, 12, 'sp4_h_r_35')
// (15, 12, 'sp4_r_v_b_17')
// (15, 13, 'sp4_h_r_47')
// (15, 13, 'sp4_r_v_b_4')
// (15, 14, 'sp4_h_r_44')
// (15, 14, 'sp4_r_v_b_38')
// (15, 15, 'local_g2_7')
// (15, 15, 'lutff_0/in_3')
// (15, 15, 'sp4_r_v_b_27')
// (15, 15, 'sp4_r_v_b_39')
// (15, 16, 'sp4_r_v_b_14')
// (15, 16, 'sp4_r_v_b_26')
// (15, 17, 'local_g1_3')
// (15, 17, 'lutff_0/in_0')
// (15, 17, 'sp4_r_v_b_15')
// (15, 17, 'sp4_r_v_b_3')
// (15, 18, 'local_g1_2')
// (15, 18, 'lutff_0/in_3')
// (15, 18, 'sp4_r_v_b_2')
// (15, 19, 'local_g2_7')
// (15, 19, 'lutff_0/in_3')
// (15, 19, 'sp4_r_v_b_39')
// (15, 20, 'sp12_h_r_8')
// (15, 20, 'sp4_h_r_16')
// (15, 20, 'sp4_r_v_b_26')
// (15, 21, 'sp4_r_v_b_15')
// (15, 22, 'sp4_r_v_b_2')
// (16, 9, 'local_g3_1')
// (16, 9, 'lutff_0/in_0')
// (16, 9, 'sp4_r_v_b_41')
// (16, 9, 'sp4_v_t_41')
// (16, 10, 'sp4_r_v_b_28')
// (16, 10, 'sp4_v_b_41')
// (16, 11, 'local_g3_4')
// (16, 11, 'lutff_0/in_3')
// (16, 11, 'sp4_r_v_b_17')
// (16, 11, 'sp4_v_b_28')
// (16, 12, 'local_g2_1')
// (16, 12, 'lutff_5/in_0')
// (16, 12, 'sp4_h_r_25')
// (16, 12, 'sp4_h_r_29')
// (16, 12, 'sp4_h_r_41')
// (16, 12, 'sp4_h_r_46')
// (16, 12, 'sp4_r_v_b_4')
// (16, 12, 'sp4_v_b_17')
// (16, 13, 'sp4_h_l_47')
// (16, 13, 'sp4_h_r_6')
// (16, 13, 'sp4_v_b_4')
// (16, 13, 'sp4_v_t_38')
// (16, 14, 'sp4_h_l_44')
// (16, 14, 'sp4_h_r_5')
// (16, 14, 'sp4_v_b_38')
// (16, 14, 'sp4_v_t_39')
// (16, 15, 'sp4_v_b_27')
// (16, 15, 'sp4_v_b_39')
// (16, 16, 'local_g1_6')
// (16, 16, 'lutff_0/in_3')
// (16, 16, 'sp4_v_b_14')
// (16, 16, 'sp4_v_b_26')
// (16, 17, 'local_g0_3')
// (16, 17, 'lutff_0/in_3')
// (16, 17, 'sp4_v_b_15')
// (16, 17, 'sp4_v_b_3')
// (16, 18, 'local_g1_2')
// (16, 18, 'lutff_0/in_3')
// (16, 18, 'sp4_v_b_2')
// (16, 18, 'sp4_v_t_39')
// (16, 19, 'local_g2_7')
// (16, 19, 'lutff_6/in_3')
// (16, 19, 'sp4_v_b_39')
// (16, 20, 'sp12_h_r_11')
// (16, 20, 'sp4_h_r_29')
// (16, 20, 'sp4_v_b_26')
// (16, 21, 'local_g0_7')
// (16, 21, 'lutff_6/in_3')
// (16, 21, 'sp4_v_b_15')
// (16, 22, 'sp4_v_b_2')
// (17, 8, 'sp4_v_t_41')
// (17, 9, 'sp4_r_v_b_40')
// (17, 9, 'sp4_v_b_41')
// (17, 10, 'sp4_r_v_b_29')
// (17, 10, 'sp4_v_b_28')
// (17, 11, 'sp4_r_v_b_16')
// (17, 11, 'sp4_v_b_17')
// (17, 12, 'sp4_h_l_41')
// (17, 12, 'sp4_h_l_46')
// (17, 12, 'sp4_h_r_36')
// (17, 12, 'sp4_h_r_40')
// (17, 12, 'sp4_h_r_7')
// (17, 12, 'sp4_r_v_b_5')
// (17, 12, 'sp4_v_b_4')
// (17, 13, 'sp4_h_r_19')
// (17, 13, 'sp4_r_v_b_36')
// (17, 14, 'sp4_h_r_16')
// (17, 14, 'sp4_r_v_b_25')
// (17, 15, 'sp4_r_v_b_12')
// (17, 16, 'sp4_r_v_b_1')
// (17, 20, 'sp12_h_r_12')
// (17, 20, 'sp4_h_r_40')
// (18, 8, 'sp4_v_t_40')
// (18, 9, 'sp4_v_b_40')
// (18, 10, 'sp4_v_b_29')
// (18, 11, 'local_g1_0')
// (18, 11, 'lutff_0/in_3')
// (18, 11, 'sp4_v_b_16')
// (18, 12, 'local_g1_2')
// (18, 12, 'lutff_0/in_3')
// (18, 12, 'sp4_h_l_36')
// (18, 12, 'sp4_h_l_40')
// (18, 12, 'sp4_h_r_18')
// (18, 12, 'sp4_v_b_5')
// (18, 12, 'sp4_v_t_36')
// (18, 13, 'sp4_h_r_30')
// (18, 13, 'sp4_v_b_36')
// (18, 14, 'sp4_h_r_29')
// (18, 14, 'sp4_v_b_25')
// (18, 15, 'local_g1_4')
// (18, 15, 'lutff_1/in_0')
// (18, 15, 'sp4_v_b_12')
// (18, 16, 'sp4_v_b_1')
// (18, 20, 'sp12_h_r_15')
// (18, 20, 'sp4_h_l_40')
// (18, 20, 'sp4_h_r_9')
// (19, 10, 'local_g2_5')
// (19, 10, 'lutff_0/in_3')
// (19, 10, 'sp4_r_v_b_37')
// (19, 11, 'local_g3_6')
// (19, 11, 'lutff_0/in_3')
// (19, 11, 'sp4_r_v_b_24')
// (19, 11, 'sp4_r_v_b_46')
// (19, 12, 'sp4_h_r_31')
// (19, 12, 'sp4_r_v_b_13')
// (19, 12, 'sp4_r_v_b_35')
// (19, 13, 'local_g2_3')
// (19, 13, 'lutff_0/in_3')
// (19, 13, 'sp4_h_r_43')
// (19, 13, 'sp4_r_v_b_0')
// (19, 13, 'sp4_r_v_b_22')
// (19, 14, 'sp4_h_r_40')
// (19, 14, 'sp4_r_v_b_11')
// (19, 15, 'local_g3_7')
// (19, 15, 'lutff_0/in_0')
// (19, 15, 'sp4_r_v_b_47')
// (19, 16, 'local_g0_1')
// (19, 16, 'lutff_0/in_1')
// (19, 16, 'sp4_r_v_b_34')
// (19, 17, 'sp4_r_v_b_23')
// (19, 18, 'sp4_r_v_b_10')
// (19, 19, 'local_g3_7')
// (19, 19, 'lutff_0/in_0')
// (19, 19, 'sp4_r_v_b_47')
// (19, 20, 'sp12_h_r_16')
// (19, 20, 'sp4_h_r_20')
// (19, 20, 'sp4_r_v_b_34')
// (19, 21, 'sp4_r_v_b_23')
// (19, 22, 'sp4_r_v_b_10')
// (19, 23, 'sp4_r_v_b_47')
// (19, 24, 'sp4_r_v_b_34')
// (19, 25, 'local_g3_7')
// (19, 25, 'lutff_0/in_0')
// (19, 25, 'sp4_r_v_b_23')
// (19, 26, 'sp4_r_v_b_10')
// (20, 9, 'sp4_r_v_b_42')
// (20, 9, 'sp4_v_t_37')
// (20, 10, 'sp4_r_v_b_31')
// (20, 10, 'sp4_v_b_37')
// (20, 10, 'sp4_v_t_46')
// (20, 11, 'sp4_r_v_b_18')
// (20, 11, 'sp4_v_b_24')
// (20, 11, 'sp4_v_b_46')
// (20, 12, 'local_g3_2')
// (20, 12, 'lutff_0/in_3')
// (20, 12, 'sp4_h_r_42')
// (20, 12, 'sp4_r_v_b_7')
// (20, 12, 'sp4_v_b_13')
// (20, 12, 'sp4_v_b_35')
// (20, 13, 'sp4_h_l_43')
// (20, 13, 'sp4_v_b_0')
// (20, 13, 'sp4_v_b_22')
// (20, 14, 'sp4_h_l_40')
// (20, 14, 'sp4_h_r_1')
// (20, 14, 'sp4_v_b_11')
// (20, 14, 'sp4_v_t_47')
// (20, 15, 'sp4_v_b_47')
// (20, 16, 'local_g3_2')
// (20, 16, 'lutff_0/in_3')
// (20, 16, 'sp4_v_b_34')
// (20, 17, 'local_g1_7')
// (20, 17, 'lutff_1/in_3')
// (20, 17, 'sp4_v_b_23')
// (20, 18, 'local_g1_2')
// (20, 18, 'lutff_1/in_0')
// (20, 18, 'lutff_2/in_1')
// (20, 18, 'sp4_v_b_10')
// (20, 18, 'sp4_v_t_47')
// (20, 19, 'local_g2_7')
// (20, 19, 'lutff_0/in_3')
// (20, 19, 'sp4_v_b_47')
// (20, 20, 'local_g0_3')
// (20, 20, 'lutff_0/in_3')
// (20, 20, 'sp12_h_r_19')
// (20, 20, 'sp4_h_r_33')
// (20, 20, 'sp4_v_b_34')
// (20, 21, 'sp4_v_b_23')
// (20, 22, 'sp4_v_b_10')
// (20, 22, 'sp4_v_t_47')
// (20, 23, 'local_g2_7')
// (20, 23, 'lutff_2/in_3')
// (20, 23, 'sp4_v_b_47')
// (20, 24, 'sp4_v_b_34')
// (20, 25, 'local_g0_7')
// (20, 25, 'lutff_0/in_3')
// (20, 25, 'sp4_v_b_23')
// (20, 26, 'sp4_v_b_10')
// (21, 8, 'sp4_v_t_42')
// (21, 9, 'sp4_v_b_42')
// (21, 10, 'sp4_v_b_31')
// (21, 11, 'local_g1_2')
// (21, 11, 'lutff_0/in_3')
// (21, 11, 'sp4_v_b_18')
// (21, 12, 'local_g1_7')
// (21, 12, 'lutff_0/in_0')
// (21, 12, 'sp4_h_l_42')
// (21, 12, 'sp4_h_r_7')
// (21, 12, 'sp4_v_b_7')
// (21, 14, 'local_g1_4')
// (21, 14, 'lutff_2/in_3')
// (21, 14, 'sp4_h_r_12')
// (21, 20, 'local_g1_4')
// (21, 20, 'lutff_0/in_3')
// (21, 20, 'sp12_h_r_20')
// (21, 20, 'sp4_h_r_44')
// (21, 21, 'sp4_r_v_b_39')
// (21, 22, 'sp4_r_v_b_26')
// (21, 23, 'sp4_r_v_b_15')
// (21, 24, 'sp4_r_v_b_2')
// (22, 12, 'local_g1_2')
// (22, 12, 'lutff_0/in_3')
// (22, 12, 'sp4_h_r_18')
// (22, 14, 'local_g2_1')
// (22, 14, 'lutff_0/in_3')
// (22, 14, 'sp4_h_r_25')
// (22, 20, 'sp12_h_r_23')
// (22, 20, 'sp4_h_l_44')
// (22, 20, 'sp4_v_t_39')
// (22, 21, 'local_g2_7')
// (22, 21, 'lutff_0/in_3')
// (22, 21, 'sp4_v_b_39')
// (22, 22, 'sp4_v_b_26')
// (22, 23, 'local_g0_7')
// (22, 23, 'lutff_0/in_3')
// (22, 23, 'sp4_v_b_15')
// (22, 24, 'sp4_v_b_2')
// (23, 8, 'sp12_v_t_23')
// (23, 9, 'sp12_v_b_23')
// (23, 10, 'sp12_v_b_20')
// (23, 11, 'sp12_v_b_19')
// (23, 12, 'local_g2_7')
// (23, 12, 'lutff_0/in_3')
// (23, 12, 'sp12_v_b_16')
// (23, 12, 'sp4_h_r_31')
// (23, 13, 'sp12_v_b_15')
// (23, 14, 'local_g3_4')
// (23, 14, 'lutff_0/in_3')
// (23, 14, 'sp12_v_b_12')
// (23, 14, 'sp4_h_r_36')
// (23, 15, 'local_g2_3')
// (23, 15, 'lutff_0/in_3')
// (23, 15, 'sp12_v_b_11')
// (23, 15, 'sp4_r_v_b_43')
// (23, 16, 'local_g1_6')
// (23, 16, 'lutff_0/in_3')
// (23, 16, 'sp12_v_b_8')
// (23, 16, 'sp4_r_v_b_30')
// (23, 17, 'sp12_v_b_7')
// (23, 17, 'sp4_r_v_b_19')
// (23, 18, 'local_g1_6')
// (23, 18, 'lutff_0/in_3')
// (23, 18, 'sp12_v_b_4')
// (23, 18, 'sp4_r_v_b_6')
// (23, 19, 'sp12_v_b_3')
// (23, 20, 'local_g3_0')
// (23, 20, 'lutff_0/in_3')
// (23, 20, 'sp12_h_l_23')
// (23, 20, 'sp12_v_b_0')
// (24, 12, 'sp4_h_r_42')
// (24, 14, 'local_g1_4')
// (24, 14, 'lutff_0/in_3')
// (24, 14, 'sp4_h_l_36')
// (24, 14, 'sp4_h_r_4')
// (24, 14, 'sp4_v_t_43')
// (24, 15, 'local_g2_3')
// (24, 15, 'lutff_0/in_3')
// (24, 15, 'sp4_v_b_43')
// (24, 16, 'sp4_v_b_30')
// (24, 17, 'local_g0_3')
// (24, 17, 'lutff_0/in_3')
// (24, 17, 'sp4_v_b_19')
// (24, 18, 'sp4_v_b_6')
// (25, 12, 'sp4_h_l_42')
// (25, 14, 'sp4_h_r_17')
// (26, 14, 'sp4_h_r_28')
// (27, 14, 'sp4_h_r_41')
// (28, 14, 'sp4_h_l_41')

wire n160;
// (8, 14, 'neigh_op_tnr_0')
// (8, 15, 'neigh_op_rgt_0')
// (8, 16, 'neigh_op_bnr_0')
// (9, 14, 'local_g1_0')
// (9, 14, 'lutff_2/in_3')
// (9, 14, 'neigh_op_top_0')
// (9, 15, 'lutff_0/out')
// (9, 16, 'neigh_op_bot_0')
// (10, 14, 'neigh_op_tnl_0')
// (10, 15, 'neigh_op_lft_0')
// (10, 16, 'neigh_op_bnl_0')

wire n161;
// (8, 14, 'neigh_op_tnr_1')
// (8, 15, 'neigh_op_rgt_1')
// (8, 16, 'neigh_op_bnr_1')
// (9, 14, 'local_g1_1')
// (9, 14, 'lutff_2/in_0')
// (9, 14, 'neigh_op_top_1')
// (9, 15, 'lutff_1/out')
// (9, 16, 'neigh_op_bot_1')
// (10, 14, 'neigh_op_tnl_1')
// (10, 15, 'neigh_op_lft_1')
// (10, 16, 'neigh_op_bnl_1')

wire n162;
// (8, 14, 'neigh_op_tnr_4')
// (8, 15, 'neigh_op_rgt_4')
// (8, 16, 'neigh_op_bnr_4')
// (9, 14, 'neigh_op_top_4')
// (9, 15, 'local_g1_4')
// (9, 15, 'lutff_0/in_3')
// (9, 15, 'lutff_4/out')
// (9, 16, 'neigh_op_bot_4')
// (10, 14, 'neigh_op_tnl_4')
// (10, 15, 'neigh_op_lft_4')
// (10, 16, 'neigh_op_bnl_4')

wire n163;
// (8, 14, 'neigh_op_tnr_6')
// (8, 15, 'neigh_op_rgt_6')
// (8, 15, 'sp4_r_v_b_44')
// (8, 16, 'neigh_op_bnr_6')
// (8, 16, 'sp4_r_v_b_33')
// (8, 17, 'sp4_r_v_b_20')
// (8, 18, 'sp4_r_v_b_9')
// (9, 14, 'neigh_op_top_6')
// (9, 14, 'sp4_h_r_2')
// (9, 14, 'sp4_v_t_44')
// (9, 15, 'lutff_6/out')
// (9, 15, 'sp4_v_b_44')
// (9, 16, 'neigh_op_bot_6')
// (9, 16, 'sp4_v_b_33')
// (9, 17, 'sp4_v_b_20')
// (9, 18, 'sp4_v_b_9')
// (10, 14, 'neigh_op_tnl_6')
// (10, 14, 'sp4_h_r_15')
// (10, 15, 'neigh_op_lft_6')
// (10, 16, 'neigh_op_bnl_6')
// (11, 14, 'sp4_h_r_26')
// (12, 14, 'sp4_h_r_39')
// (13, 14, 'sp4_h_l_39')
// (13, 14, 'sp4_h_r_2')
// (14, 14, 'sp4_h_r_15')
// (15, 14, 'local_g2_2')
// (15, 14, 'lutff_5/in_1')
// (15, 14, 'sp4_h_r_26')
// (16, 14, 'sp4_h_r_39')
// (17, 14, 'sp4_h_l_39')

wire n164;
// (8, 14, 'neigh_op_tnr_7')
// (8, 15, 'neigh_op_rgt_7')
// (8, 16, 'neigh_op_bnr_7')
// (9, 14, 'neigh_op_top_7')
// (9, 15, 'local_g2_7')
// (9, 15, 'lutff_0/in_1')
// (9, 15, 'lutff_7/out')
// (9, 16, 'neigh_op_bot_7')
// (10, 14, 'neigh_op_tnl_7')
// (10, 15, 'neigh_op_lft_7')
// (10, 16, 'neigh_op_bnl_7')

wire n165;
// (8, 14, 'sp4_r_v_b_42')
// (8, 15, 'neigh_op_tnr_1')
// (8, 15, 'sp4_r_v_b_31')
// (8, 16, 'neigh_op_rgt_1')
// (8, 16, 'sp4_r_v_b_18')
// (8, 17, 'neigh_op_bnr_1')
// (8, 17, 'sp4_r_v_b_7')
// (9, 13, 'sp4_v_t_42')
// (9, 14, 'local_g3_2')
// (9, 14, 'lutff_2/in_1')
// (9, 14, 'sp4_v_b_42')
// (9, 15, 'neigh_op_top_1')
// (9, 15, 'sp4_v_b_31')
// (9, 16, 'lutff_1/out')
// (9, 16, 'sp4_v_b_18')
// (9, 17, 'neigh_op_bot_1')
// (9, 17, 'sp4_v_b_7')
// (10, 15, 'neigh_op_tnl_1')
// (10, 16, 'neigh_op_lft_1')
// (10, 17, 'neigh_op_bnl_1')

wire n166;
// (8, 15, 'neigh_op_tnr_0')
// (8, 16, 'neigh_op_rgt_0')
// (8, 17, 'neigh_op_bnr_0')
// (9, 15, 'local_g0_0')
// (9, 15, 'lutff_0/in_0')
// (9, 15, 'neigh_op_top_0')
// (9, 16, 'lutff_0/out')
// (9, 17, 'neigh_op_bot_0')
// (10, 15, 'neigh_op_tnl_0')
// (10, 16, 'neigh_op_lft_0')
// (10, 17, 'neigh_op_bnl_0')

wire n167;
// (8, 15, 'neigh_op_tnr_2')
// (8, 16, 'neigh_op_rgt_2')
// (8, 17, 'neigh_op_bnr_2')
// (9, 15, 'local_g0_2')
// (9, 15, 'lutff_0/in_2')
// (9, 15, 'neigh_op_top_2')
// (9, 16, 'lutff_2/out')
// (9, 17, 'neigh_op_bot_2')
// (10, 15, 'neigh_op_tnl_2')
// (10, 16, 'neigh_op_lft_2')
// (10, 17, 'neigh_op_bnl_2')

wire n168;
// (8, 15, 'neigh_op_tnr_3')
// (8, 16, 'neigh_op_rgt_3')
// (8, 16, 'sp4_h_r_11')
// (8, 17, 'neigh_op_bnr_3')
// (9, 15, 'neigh_op_top_3')
// (9, 16, 'lutff_3/out')
// (9, 16, 'sp4_h_r_22')
// (9, 17, 'neigh_op_bot_3')
// (10, 15, 'neigh_op_tnl_3')
// (10, 16, 'neigh_op_lft_3')
// (10, 16, 'sp4_h_r_35')
// (10, 17, 'neigh_op_bnl_3')
// (11, 16, 'local_g2_6')
// (11, 16, 'lutff_5/in_1')
// (11, 16, 'sp4_h_r_46')
// (12, 16, 'sp4_h_l_46')

wire n169;
// (8, 15, 'neigh_op_tnr_4')
// (8, 16, 'neigh_op_rgt_4')
// (8, 17, 'neigh_op_bnr_4')
// (9, 15, 'neigh_op_top_4')
// (9, 16, 'lutff_4/out')
// (9, 16, 'sp12_h_r_0')
// (9, 17, 'neigh_op_bot_4')
// (10, 15, 'neigh_op_tnl_4')
// (10, 16, 'neigh_op_lft_4')
// (10, 16, 'sp12_h_r_3')
// (10, 17, 'neigh_op_bnl_4')
// (11, 16, 'local_g0_4')
// (11, 16, 'lutff_7/in_1')
// (11, 16, 'sp12_h_r_4')
// (12, 16, 'sp12_h_r_7')
// (13, 16, 'sp12_h_r_8')
// (14, 16, 'sp12_h_r_11')
// (15, 16, 'sp12_h_r_12')
// (16, 16, 'sp12_h_r_15')
// (17, 16, 'sp12_h_r_16')
// (18, 16, 'sp12_h_r_19')
// (19, 16, 'sp12_h_r_20')
// (20, 16, 'sp12_h_r_23')
// (21, 16, 'sp12_h_l_23')

wire n170;
// (8, 15, 'neigh_op_tnr_7')
// (8, 16, 'neigh_op_rgt_7')
// (8, 17, 'neigh_op_bnr_7')
// (9, 15, 'local_g0_7')
// (9, 15, 'lutff_6/in_3')
// (9, 15, 'neigh_op_top_7')
// (9, 16, 'lutff_7/out')
// (9, 17, 'neigh_op_bot_7')
// (10, 15, 'neigh_op_tnl_7')
// (10, 16, 'neigh_op_lft_7')
// (10, 17, 'neigh_op_bnl_7')

reg n171 = 0;
// (8, 15, 'sp12_h_r_0')
// (9, 15, 'sp12_h_r_3')
// (10, 15, 'sp12_h_r_4')
// (11, 15, 'sp12_h_r_7')
// (12, 15, 'sp12_h_r_8')
// (13, 15, 'sp12_h_r_11')
// (14, 15, 'sp12_h_r_12')
// (15, 15, 'sp12_h_r_15')
// (16, 15, 'sp12_h_r_16')
// (17, 15, 'local_g1_3')
// (17, 15, 'lutff_5/in_3')
// (17, 15, 'sp12_h_r_19')
// (18, 15, 'sp12_h_r_20')
// (19, 15, 'sp12_h_r_23')
// (20, 15, 'sp12_h_l_23')
// (20, 15, 'sp12_h_r_0')
// (21, 15, 'sp12_h_r_3')
// (22, 15, 'sp12_h_r_4')
// (23, 14, 'neigh_op_tnr_0')
// (23, 15, 'neigh_op_rgt_0')
// (23, 15, 'sp12_h_r_7')
// (23, 16, 'neigh_op_bnr_0')
// (24, 14, 'neigh_op_top_0')
// (24, 15, 'lutff_0/out')
// (24, 15, 'sp12_h_r_8')
// (24, 16, 'neigh_op_bot_0')
// (25, 14, 'neigh_op_tnl_0')
// (25, 15, 'neigh_op_lft_0')
// (25, 15, 'sp12_h_r_11')
// (25, 16, 'neigh_op_bnl_0')
// (26, 15, 'sp12_h_r_12')
// (27, 15, 'sp12_h_r_15')
// (28, 15, 'sp12_h_r_16')
// (29, 15, 'sp12_h_r_19')
// (30, 15, 'sp12_h_r_20')
// (31, 15, 'sp12_h_r_23')
// (32, 15, 'sp12_h_l_23')

wire n172;
// (8, 15, 'sp4_r_v_b_40')
// (8, 16, 'neigh_op_tnr_0')
// (8, 16, 'sp4_r_v_b_29')
// (8, 17, 'neigh_op_rgt_0')
// (8, 17, 'sp4_r_v_b_16')
// (8, 18, 'neigh_op_bnr_0')
// (8, 18, 'sp4_r_v_b_5')
// (9, 14, 'sp4_v_t_40')
// (9, 15, 'sp4_v_b_40')
// (9, 16, 'neigh_op_top_0')
// (9, 16, 'sp4_r_v_b_44')
// (9, 16, 'sp4_v_b_29')
// (9, 17, 'local_g0_2')
// (9, 17, 'lutff_0/out')
// (9, 17, 'lutff_global/cen')
// (9, 17, 'sp4_r_v_b_33')
// (9, 17, 'sp4_v_b_16')
// (9, 18, 'local_g1_3')
// (9, 18, 'lutff_global/cen')
// (9, 18, 'neigh_op_bot_0')
// (9, 18, 'sp4_h_r_11')
// (9, 18, 'sp4_r_v_b_20')
// (9, 18, 'sp4_v_b_5')
// (9, 19, 'sp4_r_v_b_9')
// (10, 15, 'sp4_v_t_44')
// (10, 16, 'neigh_op_tnl_0')
// (10, 16, 'sp4_v_b_44')
// (10, 17, 'neigh_op_lft_0')
// (10, 17, 'sp4_v_b_33')
// (10, 18, 'neigh_op_bnl_0')
// (10, 18, 'sp4_h_r_22')
// (10, 18, 'sp4_v_b_20')
// (10, 19, 'sp4_v_b_9')
// (11, 18, 'sp4_h_r_35')
// (12, 18, 'sp4_h_r_46')
// (13, 18, 'sp4_h_l_46')

reg n173 = 0;
// (8, 16, 'neigh_op_tnr_1')
// (8, 17, 'neigh_op_rgt_1')
// (8, 18, 'neigh_op_bnr_1')
// (9, 16, 'neigh_op_top_1')
// (9, 17, 'lutff_1/out')
// (9, 17, 'sp4_h_r_2')
// (9, 18, 'neigh_op_bot_1')
// (10, 16, 'neigh_op_tnl_1')
// (10, 17, 'neigh_op_lft_1')
// (10, 17, 'sp4_h_r_15')
// (10, 18, 'neigh_op_bnl_1')
// (11, 17, 'sp4_h_r_26')
// (12, 17, 'sp4_h_r_39')
// (12, 18, 'sp4_r_v_b_39')
// (12, 19, 'sp4_r_v_b_26')
// (12, 20, 'sp4_r_v_b_15')
// (12, 21, 'sp4_r_v_b_2')
// (13, 17, 'sp4_h_l_39')
// (13, 17, 'sp4_v_t_39')
// (13, 18, 'local_g2_7')
// (13, 18, 'lutff_0/in_1')
// (13, 18, 'sp4_v_b_39')
// (13, 19, 'sp4_v_b_26')
// (13, 20, 'sp4_v_b_15')
// (13, 21, 'sp4_v_b_2')

reg n174 = 0;
// (8, 16, 'neigh_op_tnr_5')
// (8, 17, 'neigh_op_rgt_5')
// (8, 17, 'sp4_r_v_b_42')
// (8, 18, 'neigh_op_bnr_5')
// (8, 18, 'sp4_r_v_b_31')
// (8, 19, 'sp4_r_v_b_18')
// (8, 20, 'sp4_r_v_b_7')
// (9, 16, 'neigh_op_top_5')
// (9, 16, 'sp4_h_r_0')
// (9, 16, 'sp4_v_t_42')
// (9, 17, 'lutff_5/out')
// (9, 17, 'sp4_v_b_42')
// (9, 18, 'neigh_op_bot_5')
// (9, 18, 'sp4_v_b_31')
// (9, 19, 'sp4_v_b_18')
// (9, 20, 'sp4_v_b_7')
// (10, 16, 'neigh_op_tnl_5')
// (10, 16, 'sp4_h_r_13')
// (10, 17, 'neigh_op_lft_5')
// (10, 18, 'neigh_op_bnl_5')
// (11, 16, 'sp4_h_r_24')
// (12, 16, 'sp4_h_r_37')
// (12, 17, 'sp4_r_v_b_37')
// (12, 18, 'sp4_r_v_b_24')
// (12, 19, 'sp4_r_v_b_13')
// (12, 20, 'sp4_r_v_b_0')
// (13, 16, 'sp4_h_l_37')
// (13, 16, 'sp4_v_t_37')
// (13, 17, 'sp4_v_b_37')
// (13, 18, 'local_g2_0')
// (13, 18, 'lutff_1/in_1')
// (13, 18, 'sp4_v_b_24')
// (13, 19, 'sp4_v_b_13')
// (13, 20, 'sp4_v_b_0')

reg n175 = 0;
// (8, 16, 'neigh_op_tnr_7')
// (8, 17, 'neigh_op_rgt_7')
// (8, 17, 'sp4_r_v_b_46')
// (8, 18, 'neigh_op_bnr_7')
// (8, 18, 'sp4_r_v_b_35')
// (8, 19, 'sp4_r_v_b_22')
// (8, 20, 'sp4_r_v_b_11')
// (9, 16, 'neigh_op_top_7')
// (9, 16, 'sp4_h_r_4')
// (9, 16, 'sp4_v_t_46')
// (9, 17, 'lutff_7/out')
// (9, 17, 'sp4_v_b_46')
// (9, 18, 'neigh_op_bot_7')
// (9, 18, 'sp4_v_b_35')
// (9, 19, 'sp4_v_b_22')
// (9, 20, 'sp4_v_b_11')
// (10, 16, 'neigh_op_tnl_7')
// (10, 16, 'sp4_h_r_17')
// (10, 17, 'neigh_op_lft_7')
// (10, 18, 'neigh_op_bnl_7')
// (11, 16, 'sp4_h_r_28')
// (12, 16, 'sp4_h_r_41')
// (12, 17, 'sp4_r_v_b_41')
// (12, 18, 'sp4_r_v_b_28')
// (12, 19, 'sp4_r_v_b_17')
// (12, 20, 'sp4_r_v_b_4')
// (13, 16, 'sp4_h_l_41')
// (13, 16, 'sp4_v_t_41')
// (13, 17, 'sp4_v_b_41')
// (13, 18, 'local_g2_4')
// (13, 18, 'lutff_3/in_1')
// (13, 18, 'sp4_v_b_28')
// (13, 19, 'sp4_v_b_17')
// (13, 20, 'sp4_v_b_4')

reg n176 = 0;
// (8, 17, 'neigh_op_tnr_0')
// (8, 18, 'neigh_op_rgt_0')
// (8, 19, 'neigh_op_bnr_0')
// (9, 17, 'neigh_op_top_0')
// (9, 18, 'lutff_0/out')
// (9, 18, 'sp4_h_r_0')
// (9, 19, 'neigh_op_bot_0')
// (10, 17, 'neigh_op_tnl_0')
// (10, 18, 'neigh_op_lft_0')
// (10, 18, 'sp4_h_r_13')
// (10, 19, 'neigh_op_bnl_0')
// (11, 18, 'sp4_h_r_24')
// (12, 18, 'sp4_h_r_37')
// (13, 18, 'local_g0_3')
// (13, 18, 'lutff_4/in_1')
// (13, 18, 'sp4_h_l_37')
// (13, 18, 'sp4_h_r_3')
// (14, 18, 'sp4_h_r_14')
// (15, 18, 'sp4_h_r_27')
// (16, 18, 'sp4_h_r_38')
// (17, 18, 'sp4_h_l_38')

reg n177 = 0;
// (8, 17, 'neigh_op_tnr_1')
// (8, 18, 'neigh_op_rgt_1')
// (8, 19, 'neigh_op_bnr_1')
// (9, 17, 'neigh_op_top_1')
// (9, 18, 'lutff_1/out')
// (9, 18, 'sp4_h_r_2')
// (9, 19, 'neigh_op_bot_1')
// (10, 17, 'neigh_op_tnl_1')
// (10, 18, 'neigh_op_lft_1')
// (10, 18, 'sp4_h_r_15')
// (10, 19, 'neigh_op_bnl_1')
// (11, 18, 'sp4_h_r_26')
// (12, 18, 'sp4_h_r_39')
// (13, 18, 'local_g0_2')
// (13, 18, 'lutff_5/in_1')
// (13, 18, 'sp4_h_l_39')
// (13, 18, 'sp4_h_r_2')
// (14, 18, 'sp4_h_r_15')
// (15, 18, 'sp4_h_r_26')
// (16, 18, 'sp4_h_r_39')
// (17, 18, 'sp4_h_l_39')

reg n178 = 0;
// (8, 17, 'neigh_op_tnr_3')
// (8, 18, 'neigh_op_rgt_3')
// (8, 18, 'sp4_h_r_11')
// (8, 19, 'neigh_op_bnr_3')
// (9, 17, 'neigh_op_top_3')
// (9, 18, 'lutff_3/out')
// (9, 18, 'sp4_h_r_22')
// (9, 19, 'neigh_op_bot_3')
// (10, 17, 'neigh_op_tnl_3')
// (10, 18, 'neigh_op_lft_3')
// (10, 18, 'sp4_h_r_35')
// (10, 19, 'neigh_op_bnl_3')
// (11, 18, 'sp4_h_r_46')
// (12, 18, 'sp4_h_l_46')
// (12, 18, 'sp4_h_r_11')
// (13, 18, 'local_g0_6')
// (13, 18, 'lutff_7/in_1')
// (13, 18, 'sp4_h_r_22')
// (14, 18, 'sp4_h_r_35')
// (15, 18, 'sp4_h_r_46')
// (16, 18, 'sp4_h_l_46')

wire n179;
// (8, 17, 'sp4_h_r_5')
// (9, 17, 'sp4_h_r_16')
// (10, 17, 'sp4_h_r_29')
// (11, 17, 'local_g2_0')
// (11, 17, 'lutff_7/in_1')
// (11, 17, 'sp4_h_r_40')
// (12, 16, 'neigh_op_tnr_0')
// (12, 17, 'neigh_op_rgt_0')
// (12, 17, 'sp4_h_l_40')
// (12, 17, 'sp4_h_r_5')
// (12, 18, 'neigh_op_bnr_0')
// (13, 13, 'sp12_v_t_23')
// (13, 14, 'sp12_v_b_23')
// (13, 15, 'sp12_v_b_20')
// (13, 16, 'neigh_op_top_0')
// (13, 16, 'sp12_v_b_19')
// (13, 17, 'lutff_0/out')
// (13, 17, 'sp12_v_b_16')
// (13, 17, 'sp4_h_r_16')
// (13, 18, 'neigh_op_bot_0')
// (13, 18, 'sp12_v_b_15')
// (13, 19, 'sp12_v_b_12')
// (13, 20, 'sp12_v_b_11')
// (13, 21, 'local_g3_0')
// (13, 21, 'lutff_3/in_2')
// (13, 21, 'sp12_v_b_8')
// (13, 22, 'sp12_v_b_7')
// (13, 23, 'sp12_v_b_4')
// (13, 24, 'sp12_v_b_3')
// (13, 25, 'sp12_v_b_0')
// (14, 16, 'neigh_op_tnl_0')
// (14, 17, 'neigh_op_lft_0')
// (14, 17, 'sp4_h_r_29')
// (14, 18, 'neigh_op_bnl_0')
// (15, 17, 'sp4_h_r_40')
// (16, 17, 'sp4_h_l_40')

reg n180 = 0;
// (8, 17, 'sp4_h_r_9')
// (9, 17, 'local_g0_4')
// (9, 17, 'lutff_0/in_0')
// (9, 17, 'sp4_h_r_20')
// (10, 17, 'sp4_h_r_33')
// (11, 17, 'sp4_h_r_44')
// (12, 17, 'sp4_h_l_44')
// (12, 17, 'sp4_h_r_1')
// (13, 17, 'sp4_h_r_12')
// (14, 17, 'sp4_h_r_25')
// (15, 10, 'sp4_r_v_b_39')
// (15, 11, 'sp4_r_v_b_26')
// (15, 12, 'neigh_op_tnr_1')
// (15, 12, 'sp4_r_v_b_15')
// (15, 13, 'neigh_op_rgt_1')
// (15, 13, 'sp4_h_r_7')
// (15, 13, 'sp4_r_v_b_2')
// (15, 14, 'neigh_op_bnr_1')
// (15, 14, 'sp4_r_v_b_45')
// (15, 15, 'sp4_r_v_b_32')
// (15, 16, 'local_g3_5')
// (15, 16, 'lutff_4/in_2')
// (15, 16, 'lutff_5/in_1')
// (15, 16, 'lutff_7/in_3')
// (15, 16, 'sp4_r_v_b_21')
// (15, 17, 'sp4_h_r_36')
// (15, 17, 'sp4_r_v_b_8')
// (16, 9, 'sp4_v_t_39')
// (16, 10, 'sp12_v_t_22')
// (16, 10, 'sp4_v_b_39')
// (16, 11, 'sp12_v_b_22')
// (16, 11, 'sp4_v_b_26')
// (16, 12, 'local_g1_1')
// (16, 12, 'lutff_0/in_0')
// (16, 12, 'lutff_7/in_1')
// (16, 12, 'neigh_op_top_1')
// (16, 12, 'sp12_v_b_21')
// (16, 12, 'sp4_v_b_15')
// (16, 13, 'local_g3_1')
// (16, 13, 'lutff_0/in_0')
// (16, 13, 'lutff_1/out')
// (16, 13, 'lutff_2/in_0')
// (16, 13, 'lutff_4/in_0')
// (16, 13, 'lutff_5/in_3')
// (16, 13, 'lutff_6/in_0')
// (16, 13, 'sp12_v_b_18')
// (16, 13, 'sp4_h_r_18')
// (16, 13, 'sp4_h_r_8')
// (16, 13, 'sp4_v_b_2')
// (16, 13, 'sp4_v_t_45')
// (16, 14, 'neigh_op_bot_1')
// (16, 14, 'sp12_v_b_17')
// (16, 14, 'sp4_v_b_45')
// (16, 15, 'local_g3_6')
// (16, 15, 'lutff_6/in_1')
// (16, 15, 'sp12_v_b_14')
// (16, 15, 'sp4_v_b_32')
// (16, 16, 'sp12_v_b_13')
// (16, 16, 'sp4_v_b_21')
// (16, 17, 'sp12_v_b_10')
// (16, 17, 'sp4_h_l_36')
// (16, 17, 'sp4_v_b_8')
// (16, 18, 'sp12_v_b_9')
// (16, 19, 'sp12_v_b_6')
// (16, 20, 'sp12_v_b_5')
// (16, 21, 'sp12_v_b_2')
// (16, 22, 'sp12_v_b_1')
// (17, 12, 'neigh_op_tnl_1')
// (17, 13, 'neigh_op_lft_1')
// (17, 13, 'sp4_h_r_21')
// (17, 13, 'sp4_h_r_31')
// (17, 14, 'neigh_op_bnl_1')
// (18, 10, 'sp4_r_v_b_36')
// (18, 11, 'sp4_r_v_b_25')
// (18, 12, 'sp4_r_v_b_12')
// (18, 13, 'sp4_h_r_32')
// (18, 13, 'sp4_h_r_42')
// (18, 13, 'sp4_r_v_b_1')
// (19, 9, 'sp4_v_t_36')
// (19, 10, 'sp4_v_b_36')
// (19, 11, 'sp4_v_b_25')
// (19, 12, 'local_g0_4')
// (19, 12, 'lutff_5/in_1')
// (19, 12, 'lutff_7/in_3')
// (19, 12, 'sp4_v_b_12')
// (19, 13, 'sp4_h_l_42')
// (19, 13, 'sp4_h_r_45')
// (19, 13, 'sp4_v_b_1')
// (19, 14, 'sp4_r_v_b_45')
// (19, 15, 'sp4_r_v_b_32')
// (19, 16, 'sp4_r_v_b_21')
// (19, 17, 'sp4_r_v_b_8')
// (20, 13, 'sp4_h_l_45')
// (20, 13, 'sp4_v_t_45')
// (20, 14, 'sp4_v_b_45')
// (20, 15, 'local_g2_0')
// (20, 15, 'local_g3_0')
// (20, 15, 'lutff_0/in_3')
// (20, 15, 'lutff_1/in_2')
// (20, 15, 'lutff_2/in_1')
// (20, 15, 'lutff_3/in_1')
// (20, 15, 'lutff_4/in_1')
// (20, 15, 'lutff_6/in_1')
// (20, 15, 'sp4_v_b_32')
// (20, 16, 'sp4_v_b_21')
// (20, 17, 'sp4_v_b_8')

reg n181 = 0;
// (8, 17, 'sp4_r_v_b_47')
// (8, 18, 'sp4_r_v_b_34')
// (8, 19, 'sp4_r_v_b_23')
// (8, 20, 'sp4_r_v_b_10')
// (9, 16, 'sp4_h_r_10')
// (9, 16, 'sp4_v_t_47')
// (9, 17, 'sp4_v_b_47')
// (9, 18, 'sp4_v_b_34')
// (9, 19, 'local_g1_7')
// (9, 19, 'lutff_2/in_2')
// (9, 19, 'sp4_v_b_23')
// (9, 20, 'sp4_v_b_10')
// (10, 14, 'sp4_r_v_b_42')
// (10, 15, 'neigh_op_tnr_1')
// (10, 15, 'sp4_r_v_b_31')
// (10, 16, 'neigh_op_rgt_1')
// (10, 16, 'sp4_h_r_23')
// (10, 16, 'sp4_r_v_b_18')
// (10, 17, 'neigh_op_bnr_1')
// (10, 17, 'sp4_r_v_b_7')
// (10, 18, 'sp4_r_v_b_38')
// (10, 19, 'sp4_r_v_b_27')
// (10, 20, 'sp4_r_v_b_14')
// (10, 21, 'sp4_r_v_b_3')
// (11, 13, 'sp4_v_t_42')
// (11, 14, 'sp4_v_b_42')
// (11, 15, 'neigh_op_top_1')
// (11, 15, 'sp4_v_b_31')
// (11, 16, 'local_g0_1')
// (11, 16, 'lutff_1/in_0')
// (11, 16, 'lutff_1/out')
// (11, 16, 'sp4_h_r_34')
// (11, 16, 'sp4_v_b_18')
// (11, 17, 'neigh_op_bot_1')
// (11, 17, 'sp4_v_b_7')
// (11, 17, 'sp4_v_t_38')
// (11, 18, 'sp4_v_b_38')
// (11, 19, 'sp4_v_b_27')
// (11, 20, 'sp4_v_b_14')
// (11, 21, 'sp4_h_r_9')
// (11, 21, 'sp4_v_b_3')
// (12, 15, 'neigh_op_tnl_1')
// (12, 16, 'neigh_op_lft_1')
// (12, 16, 'sp4_h_r_47')
// (12, 17, 'neigh_op_bnl_1')
// (12, 21, 'sp4_h_r_20')
// (13, 16, 'sp4_h_l_47')
// (13, 21, 'local_g2_1')
// (13, 21, 'lutff_7/in_0')
// (13, 21, 'sp4_h_r_33')
// (14, 21, 'sp4_h_r_44')
// (15, 21, 'sp4_h_l_44')

wire n182;
// (8, 18, 'sp12_h_r_1')
// (9, 18, 'sp12_h_r_2')
// (10, 18, 'sp12_h_r_5')
// (11, 18, 'sp12_h_r_6')
// (12, 17, 'neigh_op_tnr_1')
// (12, 18, 'neigh_op_rgt_1')
// (12, 18, 'sp12_h_r_9')
// (12, 19, 'neigh_op_bnr_1')
// (13, 17, 'neigh_op_top_1')
// (13, 18, 'local_g2_1')
// (13, 18, 'lutff_1/in_2')
// (13, 18, 'lutff_1/out')
// (13, 18, 'sp12_h_r_10')
// (13, 19, 'neigh_op_bot_1')
// (14, 17, 'neigh_op_tnl_1')
// (14, 18, 'neigh_op_lft_1')
// (14, 18, 'sp12_h_r_13')
// (14, 19, 'neigh_op_bnl_1')
// (15, 18, 'sp12_h_r_14')
// (16, 18, 'sp12_h_r_17')
// (17, 18, 'local_g0_2')
// (17, 18, 'lutff_1/in_1')
// (17, 18, 'sp12_h_r_18')
// (18, 18, 'sp12_h_r_21')
// (19, 18, 'sp12_h_r_22')
// (20, 18, 'sp12_h_l_22')

reg n183 = 0;
// (8, 18, 'sp4_h_r_3')
// (9, 18, 'sp4_h_r_14')
// (10, 17, 'sp4_h_r_5')
// (10, 18, 'sp4_h_r_27')
// (11, 17, 'local_g1_0')
// (11, 17, 'lutff_6/in_3')
// (11, 17, 'sp4_h_r_16')
// (11, 18, 'local_g2_6')
// (11, 18, 'lutff_4/in_2')
// (11, 18, 'sp4_h_r_38')
// (11, 19, 'sp4_r_v_b_43')
// (11, 20, 'sp4_r_v_b_30')
// (11, 21, 'sp4_r_v_b_19')
// (11, 22, 'sp4_r_v_b_6')
// (12, 17, 'sp4_h_r_29')
// (12, 18, 'sp4_h_l_38')
// (12, 18, 'sp4_h_r_0')
// (12, 18, 'sp4_v_t_43')
// (12, 19, 'sp4_v_b_43')
// (12, 20, 'sp4_v_b_30')
// (12, 21, 'local_g1_3')
// (12, 21, 'lutff_4/in_2')
// (12, 21, 'sp4_v_b_19')
// (12, 22, 'sp4_h_r_6')
// (12, 22, 'sp4_v_b_6')
// (13, 17, 'local_g2_4')
// (13, 17, 'lutff_5/in_1')
// (13, 17, 'lutff_7/in_1')
// (13, 17, 'neigh_op_tnr_4')
// (13, 17, 'sp4_h_r_40')
// (13, 18, 'local_g3_4')
// (13, 18, 'lutff_4/in_3')
// (13, 18, 'neigh_op_rgt_4')
// (13, 18, 'sp4_h_r_13')
// (13, 18, 'sp4_r_v_b_40')
// (13, 19, 'neigh_op_bnr_4')
// (13, 19, 'sp4_r_v_b_29')
// (13, 20, 'sp4_r_v_b_16')
// (13, 21, 'local_g1_5')
// (13, 21, 'lutff_3/in_3')
// (13, 21, 'sp4_r_v_b_5')
// (13, 22, 'local_g0_3')
// (13, 22, 'lutff_4/in_1')
// (13, 22, 'sp4_h_r_19')
// (14, 17, 'neigh_op_top_4')
// (14, 17, 'sp4_h_l_40')
// (14, 17, 'sp4_v_t_40')
// (14, 18, 'local_g3_4')
// (14, 18, 'lutff_4/in_1')
// (14, 18, 'lutff_4/out')
// (14, 18, 'sp4_h_r_24')
// (14, 18, 'sp4_v_b_40')
// (14, 19, 'neigh_op_bot_4')
// (14, 19, 'sp4_v_b_29')
// (14, 20, 'sp4_v_b_16')
// (14, 21, 'sp4_v_b_5')
// (14, 22, 'sp4_h_r_30')
// (15, 17, 'neigh_op_tnl_4')
// (15, 18, 'neigh_op_lft_4')
// (15, 18, 'sp4_h_r_37')
// (15, 19, 'neigh_op_bnl_4')
// (15, 19, 'sp4_r_v_b_37')
// (15, 20, 'local_g0_0')
// (15, 20, 'lutff_4/in_2')
// (15, 20, 'sp4_r_v_b_24')
// (15, 21, 'sp4_r_v_b_13')
// (15, 22, 'sp4_h_r_43')
// (15, 22, 'sp4_r_v_b_0')
// (16, 18, 'sp4_h_l_37')
// (16, 18, 'sp4_v_t_37')
// (16, 19, 'sp4_v_b_37')
// (16, 20, 'sp4_v_b_24')
// (16, 21, 'sp4_v_b_13')
// (16, 22, 'sp4_h_l_43')
// (16, 22, 'sp4_h_r_6')
// (16, 22, 'sp4_v_b_0')
// (17, 22, 'local_g0_3')
// (17, 22, 'lutff_4/in_1')
// (17, 22, 'sp4_h_r_19')
// (18, 22, 'sp4_h_r_30')
// (19, 22, 'sp4_h_r_43')
// (20, 22, 'sp4_h_l_43')

reg n184 = 0;
// (8, 18, 'sp4_h_r_6')
// (8, 18, 'sp4_h_r_9')
// (9, 18, 'sp4_h_r_19')
// (9, 18, 'sp4_h_r_20')
// (10, 18, 'sp4_h_r_30')
// (10, 18, 'sp4_h_r_33')
// (11, 18, 'local_g2_3')
// (11, 18, 'lutff_7/in_2')
// (11, 18, 'sp4_h_r_43')
// (11, 18, 'sp4_h_r_44')
// (11, 19, 'sp4_r_v_b_39')
// (11, 20, 'sp4_r_v_b_26')
// (11, 21, 'sp4_r_v_b_15')
// (11, 22, 'sp4_r_v_b_2')
// (12, 18, 'sp4_h_l_43')
// (12, 18, 'sp4_h_l_44')
// (12, 18, 'sp4_h_r_6')
// (12, 18, 'sp4_v_t_39')
// (12, 19, 'sp4_v_b_39')
// (12, 20, 'sp4_v_b_26')
// (12, 21, 'local_g0_7')
// (12, 21, 'lutff_7/in_2')
// (12, 21, 'sp4_v_b_15')
// (12, 22, 'sp4_h_r_2')
// (12, 22, 'sp4_v_b_2')
// (13, 17, 'local_g2_7')
// (13, 17, 'local_g3_7')
// (13, 17, 'lutff_0/in_2')
// (13, 17, 'lutff_1/in_2')
// (13, 17, 'lutff_5/in_2')
// (13, 17, 'neigh_op_tnr_7')
// (13, 18, 'local_g3_7')
// (13, 18, 'lutff_7/in_3')
// (13, 18, 'neigh_op_rgt_7')
// (13, 18, 'sp4_h_r_19')
// (13, 19, 'neigh_op_bnr_7')
// (13, 22, 'local_g0_7')
// (13, 22, 'lutff_7/in_2')
// (13, 22, 'sp4_h_r_15')
// (14, 17, 'neigh_op_top_7')
// (14, 18, 'local_g3_7')
// (14, 18, 'lutff_7/in_1')
// (14, 18, 'lutff_7/out')
// (14, 18, 'sp4_h_r_30')
// (14, 19, 'neigh_op_bot_7')
// (14, 22, 'sp4_h_r_26')
// (15, 17, 'neigh_op_tnl_7')
// (15, 18, 'neigh_op_lft_7')
// (15, 18, 'sp4_h_r_43')
// (15, 19, 'neigh_op_bnl_7')
// (15, 19, 'sp4_r_v_b_46')
// (15, 20, 'local_g2_3')
// (15, 20, 'lutff_7/in_2')
// (15, 20, 'sp4_r_v_b_35')
// (15, 21, 'sp4_r_v_b_22')
// (15, 22, 'sp4_h_r_39')
// (15, 22, 'sp4_r_v_b_11')
// (16, 18, 'sp4_h_l_43')
// (16, 18, 'sp4_v_t_46')
// (16, 19, 'sp4_v_b_46')
// (16, 20, 'sp4_v_b_35')
// (16, 21, 'sp4_v_b_22')
// (16, 22, 'sp4_h_l_39')
// (16, 22, 'sp4_h_r_5')
// (16, 22, 'sp4_v_b_11')
// (17, 22, 'local_g0_0')
// (17, 22, 'lutff_7/in_1')
// (17, 22, 'sp4_h_r_16')
// (18, 22, 'sp4_h_r_29')
// (19, 22, 'sp4_h_r_40')
// (20, 22, 'sp4_h_l_40')

reg n185 = 0;
// (8, 18, 'sp4_h_r_7')
// (9, 18, 'sp4_h_r_18')
// (10, 18, 'sp4_h_r_31')
// (11, 18, 'local_g2_2')
// (11, 18, 'lutff_6/in_2')
// (11, 18, 'sp4_h_r_42')
// (11, 19, 'sp4_r_v_b_41')
// (11, 20, 'sp4_r_v_b_28')
// (11, 21, 'sp4_r_v_b_17')
// (11, 22, 'sp4_r_v_b_4')
// (12, 18, 'sp4_h_l_42')
// (12, 18, 'sp4_h_r_4')
// (12, 18, 'sp4_v_t_41')
// (12, 19, 'sp4_v_b_41')
// (12, 20, 'sp4_v_b_28')
// (12, 21, 'local_g1_1')
// (12, 21, 'lutff_6/in_2')
// (12, 21, 'sp4_v_b_17')
// (12, 22, 'sp4_h_r_4')
// (12, 22, 'sp4_v_b_4')
// (13, 17, 'local_g3_6')
// (13, 17, 'lutff_0/in_1')
// (13, 17, 'lutff_1/in_0')
// (13, 17, 'lutff_5/in_0')
// (13, 17, 'neigh_op_tnr_6')
// (13, 18, 'local_g3_6')
// (13, 18, 'lutff_6/in_3')
// (13, 18, 'neigh_op_rgt_6')
// (13, 18, 'sp4_h_r_17')
// (13, 19, 'neigh_op_bnr_6')
// (13, 22, 'local_g1_1')
// (13, 22, 'lutff_6/in_2')
// (13, 22, 'sp4_h_r_17')
// (14, 17, 'neigh_op_top_6')
// (14, 18, 'local_g1_6')
// (14, 18, 'lutff_6/in_1')
// (14, 18, 'lutff_6/out')
// (14, 18, 'sp4_h_r_28')
// (14, 19, 'neigh_op_bot_6')
// (14, 22, 'sp4_h_r_28')
// (15, 17, 'neigh_op_tnl_6')
// (15, 18, 'neigh_op_lft_6')
// (15, 18, 'sp4_h_r_41')
// (15, 19, 'neigh_op_bnl_6')
// (15, 19, 'sp4_r_v_b_44')
// (15, 20, 'local_g2_1')
// (15, 20, 'lutff_6/in_1')
// (15, 20, 'sp4_r_v_b_33')
// (15, 21, 'sp4_r_v_b_20')
// (15, 22, 'sp4_h_r_41')
// (15, 22, 'sp4_r_v_b_9')
// (16, 18, 'sp4_h_l_41')
// (16, 18, 'sp4_v_t_44')
// (16, 19, 'sp4_v_b_44')
// (16, 20, 'sp4_v_b_33')
// (16, 21, 'sp4_v_b_20')
// (16, 22, 'sp4_h_l_41')
// (16, 22, 'sp4_h_r_3')
// (16, 22, 'sp4_v_b_9')
// (17, 22, 'local_g1_6')
// (17, 22, 'lutff_6/in_1')
// (17, 22, 'sp4_h_r_14')
// (18, 22, 'sp4_h_r_27')
// (19, 22, 'sp4_h_r_38')
// (20, 22, 'sp4_h_l_38')

wire n186;
// (8, 19, 'sp12_h_r_1')
// (9, 19, 'sp12_h_r_2')
// (10, 19, 'sp12_h_r_5')
// (11, 19, 'sp12_h_r_6')
// (12, 18, 'neigh_op_tnr_1')
// (12, 19, 'neigh_op_rgt_1')
// (12, 19, 'sp12_h_r_9')
// (12, 20, 'neigh_op_bnr_1')
// (13, 18, 'neigh_op_top_1')
// (13, 19, 'local_g1_1')
// (13, 19, 'lutff_1/in_1')
// (13, 19, 'lutff_1/out')
// (13, 19, 'sp12_h_r_10')
// (13, 20, 'neigh_op_bot_1')
// (14, 18, 'neigh_op_tnl_1')
// (14, 19, 'neigh_op_lft_1')
// (14, 19, 'sp12_h_r_13')
// (14, 20, 'neigh_op_bnl_1')
// (15, 19, 'sp12_h_r_14')
// (16, 19, 'sp12_h_r_17')
// (17, 19, 'local_g0_2')
// (17, 19, 'lutff_1/in_1')
// (17, 19, 'sp12_h_r_18')
// (18, 19, 'sp12_h_r_21')
// (19, 19, 'sp12_h_r_22')
// (20, 19, 'sp12_h_l_22')

reg n187 = 0;
// (8, 19, 'sp4_h_r_3')
// (9, 19, 'sp4_h_r_14')
// (10, 19, 'sp4_h_r_27')
// (11, 19, 'local_g2_6')
// (11, 19, 'lutff_4/in_2')
// (11, 19, 'sp4_h_r_38')
// (11, 20, 'sp4_r_v_b_38')
// (11, 21, 'sp4_r_v_b_27')
// (11, 22, 'sp4_r_v_b_14')
// (11, 23, 'sp4_r_v_b_3')
// (12, 19, 'sp4_h_l_38')
// (12, 19, 'sp4_h_r_0')
// (12, 19, 'sp4_v_t_38')
// (12, 20, 'sp4_v_b_38')
// (12, 21, 'sp4_v_b_27')
// (12, 22, 'local_g0_6')
// (12, 22, 'lutff_4/in_2')
// (12, 22, 'sp4_v_b_14')
// (12, 23, 'sp4_h_r_5')
// (12, 23, 'sp4_v_b_3')
// (13, 16, 'sp4_r_v_b_45')
// (13, 17, 'sp4_r_v_b_32')
// (13, 18, 'neigh_op_tnr_4')
// (13, 18, 'sp4_r_v_b_21')
// (13, 19, 'local_g2_4')
// (13, 19, 'lutff_4/in_0')
// (13, 19, 'neigh_op_rgt_4')
// (13, 19, 'sp4_h_r_13')
// (13, 19, 'sp4_r_v_b_8')
// (13, 20, 'neigh_op_bnr_4')
// (13, 23, 'local_g0_0')
// (13, 23, 'lutff_4/in_2')
// (13, 23, 'sp4_h_r_16')
// (14, 15, 'sp4_v_t_45')
// (14, 16, 'sp4_v_b_45')
// (14, 17, 'local_g3_0')
// (14, 17, 'lutff_2/in_3')
// (14, 17, 'sp4_v_b_32')
// (14, 18, 'neigh_op_top_4')
// (14, 18, 'sp4_v_b_21')
// (14, 19, 'local_g3_4')
// (14, 19, 'lutff_4/in_1')
// (14, 19, 'lutff_4/out')
// (14, 19, 'sp4_h_r_24')
// (14, 19, 'sp4_v_b_8')
// (14, 20, 'neigh_op_bot_4')
// (14, 23, 'sp4_h_r_29')
// (15, 18, 'neigh_op_tnl_4')
// (15, 19, 'neigh_op_lft_4')
// (15, 19, 'sp4_h_r_37')
// (15, 20, 'neigh_op_bnl_4')
// (15, 20, 'sp4_r_v_b_37')
// (15, 21, 'local_g0_0')
// (15, 21, 'lutff_4/in_2')
// (15, 21, 'sp4_r_v_b_24')
// (15, 22, 'sp4_r_v_b_13')
// (15, 23, 'sp4_h_r_40')
// (15, 23, 'sp4_r_v_b_0')
// (16, 19, 'sp4_h_l_37')
// (16, 19, 'sp4_v_t_37')
// (16, 20, 'sp4_v_b_37')
// (16, 21, 'sp4_v_b_24')
// (16, 22, 'sp4_v_b_13')
// (16, 23, 'sp4_h_l_40')
// (16, 23, 'sp4_h_r_6')
// (16, 23, 'sp4_v_b_0')
// (17, 23, 'local_g0_3')
// (17, 23, 'lutff_4/in_1')
// (17, 23, 'sp4_h_r_19')
// (18, 23, 'sp4_h_r_30')
// (19, 23, 'sp4_h_r_43')
// (20, 23, 'sp4_h_l_43')

reg n188 = 0;
// (8, 19, 'sp4_h_r_7')
// (9, 19, 'sp4_h_r_18')
// (10, 19, 'sp4_h_r_31')
// (11, 19, 'local_g2_2')
// (11, 19, 'lutff_6/in_2')
// (11, 19, 'sp4_h_r_42')
// (11, 20, 'sp4_r_v_b_47')
// (11, 21, 'sp4_r_v_b_34')
// (11, 22, 'sp4_r_v_b_23')
// (11, 23, 'sp4_r_v_b_10')
// (12, 19, 'sp4_h_l_42')
// (12, 19, 'sp4_h_r_4')
// (12, 19, 'sp4_v_t_47')
// (12, 20, 'sp4_v_b_47')
// (12, 21, 'sp4_v_b_34')
// (12, 22, 'local_g1_7')
// (12, 22, 'lutff_6/in_2')
// (12, 22, 'sp4_v_b_23')
// (12, 23, 'sp4_h_r_9')
// (12, 23, 'sp4_v_b_10')
// (13, 17, 'sp4_r_v_b_36')
// (13, 18, 'neigh_op_tnr_6')
// (13, 18, 'sp4_r_v_b_25')
// (13, 19, 'local_g3_6')
// (13, 19, 'lutff_6/in_3')
// (13, 19, 'neigh_op_rgt_6')
// (13, 19, 'sp4_h_r_17')
// (13, 19, 'sp4_r_v_b_12')
// (13, 20, 'neigh_op_bnr_6')
// (13, 20, 'sp4_r_v_b_1')
// (13, 23, 'local_g0_4')
// (13, 23, 'lutff_6/in_2')
// (13, 23, 'sp4_h_r_20')
// (14, 16, 'sp4_v_t_36')
// (14, 17, 'local_g2_4')
// (14, 17, 'lutff_2/in_0')
// (14, 17, 'sp4_v_b_36')
// (14, 18, 'neigh_op_top_6')
// (14, 18, 'sp4_v_b_25')
// (14, 19, 'local_g1_6')
// (14, 19, 'lutff_6/in_1')
// (14, 19, 'lutff_6/out')
// (14, 19, 'sp4_h_r_28')
// (14, 19, 'sp4_v_b_12')
// (14, 20, 'neigh_op_bot_6')
// (14, 20, 'sp4_v_b_1')
// (14, 23, 'sp4_h_r_33')
// (15, 18, 'neigh_op_tnl_6')
// (15, 19, 'neigh_op_lft_6')
// (15, 19, 'sp4_h_r_41')
// (15, 20, 'neigh_op_bnl_6')
// (15, 20, 'sp4_r_v_b_41')
// (15, 21, 'local_g0_4')
// (15, 21, 'lutff_6/in_2')
// (15, 21, 'sp4_r_v_b_28')
// (15, 22, 'sp4_r_v_b_17')
// (15, 23, 'sp4_h_r_44')
// (15, 23, 'sp4_r_v_b_4')
// (16, 19, 'sp4_h_l_41')
// (16, 19, 'sp4_v_t_41')
// (16, 20, 'sp4_v_b_41')
// (16, 21, 'sp4_v_b_28')
// (16, 22, 'sp4_v_b_17')
// (16, 23, 'sp4_h_l_44')
// (16, 23, 'sp4_h_r_10')
// (16, 23, 'sp4_v_b_4')
// (17, 23, 'local_g0_7')
// (17, 23, 'lutff_6/in_1')
// (17, 23, 'sp4_h_r_23')
// (18, 23, 'sp4_h_r_34')
// (19, 23, 'sp4_h_r_47')
// (20, 23, 'sp4_h_l_47')

reg n189 = 0;
// (8, 20, 'sp4_h_r_3')
// (9, 20, 'sp4_h_r_14')
// (10, 20, 'sp4_h_r_27')
// (11, 20, 'local_g2_6')
// (11, 20, 'lutff_4/in_2')
// (11, 20, 'sp4_h_r_38')
// (11, 21, 'sp4_r_v_b_38')
// (11, 22, 'sp4_r_v_b_27')
// (11, 23, 'sp4_r_v_b_14')
// (11, 24, 'sp4_r_v_b_3')
// (12, 20, 'sp4_h_l_38')
// (12, 20, 'sp4_h_r_0')
// (12, 20, 'sp4_v_t_38')
// (12, 21, 'sp4_v_b_38')
// (12, 22, 'sp4_v_b_27')
// (12, 23, 'local_g0_6')
// (12, 23, 'lutff_4/in_2')
// (12, 23, 'sp4_v_b_14')
// (12, 24, 'sp4_h_r_0')
// (12, 24, 'sp4_v_b_3')
// (13, 17, 'sp4_r_v_b_45')
// (13, 18, 'sp4_r_v_b_32')
// (13, 19, 'neigh_op_tnr_4')
// (13, 19, 'sp4_r_v_b_21')
// (13, 20, 'local_g3_4')
// (13, 20, 'lutff_4/in_3')
// (13, 20, 'neigh_op_rgt_4')
// (13, 20, 'sp4_h_r_13')
// (13, 20, 'sp4_r_v_b_8')
// (13, 21, 'neigh_op_bnr_4')
// (13, 24, 'local_g1_5')
// (13, 24, 'lutff_4/in_2')
// (13, 24, 'sp4_h_r_13')
// (14, 16, 'sp4_v_t_45')
// (14, 17, 'local_g3_5')
// (14, 17, 'lutff_1/in_1')
// (14, 17, 'sp4_v_b_45')
// (14, 18, 'sp4_v_b_32')
// (14, 19, 'neigh_op_top_4')
// (14, 19, 'sp4_v_b_21')
// (14, 20, 'local_g3_4')
// (14, 20, 'lutff_4/in_1')
// (14, 20, 'lutff_4/out')
// (14, 20, 'sp4_h_r_24')
// (14, 20, 'sp4_h_r_8')
// (14, 20, 'sp4_v_b_8')
// (14, 21, 'neigh_op_bot_4')
// (14, 24, 'sp4_h_r_24')
// (15, 19, 'neigh_op_tnl_4')
// (15, 20, 'neigh_op_lft_4')
// (15, 20, 'sp4_h_r_21')
// (15, 20, 'sp4_h_r_37')
// (15, 21, 'neigh_op_bnl_4')
// (15, 21, 'sp4_r_v_b_37')
// (15, 22, 'local_g1_0')
// (15, 22, 'lutff_4/in_1')
// (15, 22, 'sp4_r_v_b_24')
// (15, 23, 'sp4_r_v_b_13')
// (15, 24, 'sp4_h_r_37')
// (15, 24, 'sp4_r_v_b_0')
// (16, 20, 'sp4_h_l_37')
// (16, 20, 'sp4_h_r_32')
// (16, 20, 'sp4_v_t_37')
// (16, 21, 'sp4_v_b_37')
// (16, 22, 'sp4_v_b_24')
// (16, 23, 'sp4_v_b_13')
// (16, 24, 'sp4_h_l_37')
// (16, 24, 'sp4_h_r_6')
// (16, 24, 'sp4_v_b_0')
// (17, 20, 'local_g3_5')
// (17, 20, 'lutff_4/in_0')
// (17, 20, 'sp4_h_r_45')
// (17, 24, 'local_g0_3')
// (17, 24, 'lutff_4/in_1')
// (17, 24, 'sp4_h_r_19')
// (18, 20, 'sp4_h_l_45')
// (18, 24, 'sp4_h_r_30')
// (19, 24, 'sp4_h_r_43')
// (20, 24, 'sp4_h_l_43')

reg n190 = 0;
// (8, 20, 'sp4_h_r_7')
// (9, 20, 'sp4_h_r_18')
// (10, 20, 'sp4_h_r_31')
// (11, 20, 'local_g2_2')
// (11, 20, 'lutff_6/in_2')
// (11, 20, 'sp4_h_r_42')
// (12, 20, 'sp12_h_r_0')
// (12, 20, 'sp12_v_t_23')
// (12, 20, 'sp4_h_l_42')
// (12, 20, 'sp4_h_r_4')
// (12, 21, 'sp12_v_b_23')
// (12, 22, 'sp12_v_b_20')
// (12, 23, 'local_g3_3')
// (12, 23, 'lutff_6/in_2')
// (12, 23, 'sp12_v_b_19')
// (12, 24, 'sp12_v_b_16')
// (12, 24, 'sp4_h_r_9')
// (12, 25, 'sp12_v_b_15')
// (12, 26, 'sp12_v_b_12')
// (12, 27, 'sp12_v_b_11')
// (12, 28, 'sp12_v_b_8')
// (12, 29, 'sp12_v_b_7')
// (12, 30, 'sp12_v_b_4')
// (12, 31, 'sp12_v_b_3')
// (12, 32, 'sp12_v_b_0')
// (13, 19, 'neigh_op_tnr_6')
// (13, 20, 'local_g2_6')
// (13, 20, 'lutff_6/in_0')
// (13, 20, 'neigh_op_rgt_6')
// (13, 20, 'sp12_h_r_3')
// (13, 20, 'sp4_h_r_17')
// (13, 21, 'neigh_op_bnr_6')
// (13, 24, 'local_g0_4')
// (13, 24, 'lutff_6/in_2')
// (13, 24, 'sp4_h_r_20')
// (14, 14, 'sp12_v_t_23')
// (14, 15, 'sp12_v_b_23')
// (14, 16, 'sp12_v_b_20')
// (14, 17, 'local_g2_3')
// (14, 17, 'lutff_1/in_2')
// (14, 17, 'sp12_v_b_19')
// (14, 18, 'sp12_v_b_16')
// (14, 19, 'neigh_op_top_6')
// (14, 19, 'sp12_v_b_15')
// (14, 20, 'local_g1_6')
// (14, 20, 'lutff_6/in_1')
// (14, 20, 'lutff_6/out')
// (14, 20, 'sp12_h_r_4')
// (14, 20, 'sp12_v_b_12')
// (14, 20, 'sp4_h_r_28')
// (14, 21, 'neigh_op_bot_6')
// (14, 21, 'sp12_v_b_11')
// (14, 22, 'sp12_v_b_8')
// (14, 23, 'sp12_v_b_7')
// (14, 24, 'sp12_v_b_4')
// (14, 24, 'sp4_h_r_33')
// (14, 25, 'sp12_v_b_3')
// (14, 26, 'sp12_v_b_0')
// (15, 19, 'neigh_op_tnl_6')
// (15, 20, 'neigh_op_lft_6')
// (15, 20, 'sp12_h_r_7')
// (15, 20, 'sp4_h_r_41')
// (15, 21, 'neigh_op_bnl_6')
// (15, 21, 'sp4_r_v_b_41')
// (15, 22, 'local_g1_4')
// (15, 22, 'lutff_6/in_1')
// (15, 22, 'sp4_r_v_b_28')
// (15, 23, 'sp4_r_v_b_17')
// (15, 24, 'sp4_h_r_44')
// (15, 24, 'sp4_r_v_b_4')
// (16, 20, 'sp12_h_r_8')
// (16, 20, 'sp4_h_l_41')
// (16, 20, 'sp4_v_t_41')
// (16, 21, 'sp4_v_b_41')
// (16, 22, 'sp4_v_b_28')
// (16, 23, 'sp4_v_b_17')
// (16, 24, 'sp4_h_l_44')
// (16, 24, 'sp4_h_r_4')
// (16, 24, 'sp4_v_b_4')
// (17, 20, 'local_g0_3')
// (17, 20, 'lutff_6/in_3')
// (17, 20, 'sp12_h_r_11')
// (17, 24, 'local_g0_1')
// (17, 24, 'lutff_6/in_1')
// (17, 24, 'sp4_h_r_17')
// (18, 20, 'sp12_h_r_12')
// (18, 24, 'sp4_h_r_28')
// (19, 20, 'sp12_h_r_15')
// (19, 24, 'sp4_h_r_41')
// (20, 20, 'sp12_h_r_16')
// (20, 24, 'sp4_h_l_41')
// (21, 20, 'sp12_h_r_19')
// (22, 20, 'sp12_h_r_20')
// (23, 20, 'sp12_h_r_23')
// (24, 20, 'sp12_h_l_23')

reg io_33_5_0 = 0;
// (8, 21, 'sp12_h_r_0')
// (9, 21, 'sp12_h_r_3')
// (10, 21, 'sp12_h_r_4')
// (11, 21, 'sp12_h_r_7')
// (12, 21, 'sp12_h_r_8')
// (13, 21, 'sp12_h_r_11')
// (14, 21, 'sp12_h_r_12')
// (15, 21, 'sp12_h_r_15')
// (16, 21, 'sp12_h_r_16')
// (17, 20, 'neigh_op_tnr_6')
// (17, 21, 'neigh_op_rgt_6')
// (17, 21, 'sp12_h_r_19')
// (17, 22, 'neigh_op_bnr_6')
// (18, 20, 'neigh_op_top_6')
// (18, 21, 'lutff_6/out')
// (18, 21, 'sp12_h_r_20')
// (18, 22, 'neigh_op_bot_6')
// (19, 20, 'neigh_op_tnl_6')
// (19, 21, 'neigh_op_lft_6')
// (19, 21, 'sp12_h_r_23')
// (19, 22, 'neigh_op_bnl_6')
// (20, 9, 'sp12_h_r_0')
// (20, 9, 'sp12_v_t_23')
// (20, 10, 'sp12_v_b_23')
// (20, 11, 'sp12_v_b_20')
// (20, 12, 'sp12_v_b_19')
// (20, 13, 'sp12_v_b_16')
// (20, 14, 'sp12_v_b_15')
// (20, 15, 'sp12_v_b_12')
// (20, 16, 'sp12_v_b_11')
// (20, 17, 'sp12_v_b_8')
// (20, 18, 'sp12_v_b_7')
// (20, 19, 'sp12_v_b_4')
// (20, 20, 'sp12_v_b_3')
// (20, 21, 'sp12_h_l_23')
// (20, 21, 'sp12_v_b_0')
// (21, 9, 'sp12_h_r_3')
// (22, 9, 'sp12_h_r_4')
// (23, 9, 'sp12_h_r_7')
// (24, 9, 'sp12_h_r_8')
// (25, 9, 'sp12_h_r_11')
// (26, 9, 'sp12_h_r_12')
// (27, 9, 'sp12_h_r_15')
// (27, 9, 'sp4_h_r_9')
// (28, 9, 'sp12_h_r_16')
// (28, 9, 'sp4_h_r_20')
// (29, 9, 'sp12_h_r_19')
// (29, 9, 'sp4_h_r_33')
// (30, 6, 'sp4_r_v_b_38')
// (30, 7, 'sp4_r_v_b_27')
// (30, 8, 'sp4_r_v_b_14')
// (30, 9, 'sp12_h_r_20')
// (30, 9, 'sp4_h_r_44')
// (30, 9, 'sp4_r_v_b_3')
// (31, 5, 'sp4_h_r_8')
// (31, 5, 'sp4_v_t_38')
// (31, 6, 'sp4_v_b_38')
// (31, 7, 'sp4_v_b_27')
// (31, 8, 'sp4_v_b_14')
// (31, 9, 'sp12_h_r_23')
// (31, 9, 'sp4_h_l_44')
// (31, 9, 'sp4_v_b_3')
// (32, 5, 'sp4_h_r_21')
// (32, 9, 'sp12_h_l_23')
// (33, 5, 'io_0/D_OUT_0')
// (33, 5, 'io_0/PAD')
// (33, 5, 'local_g1_5')
// (33, 5, 'span4_horz_21')

reg n192 = 0;
// (8, 24, 'sp12_h_r_0')
// (9, 24, 'sp12_h_r_3')
// (10, 24, 'sp12_h_r_4')
// (11, 24, 'sp12_h_r_7')
// (12, 24, 'sp12_h_r_8')
// (13, 24, 'sp12_h_r_11')
// (14, 24, 'sp12_h_r_12')
// (15, 23, 'neigh_op_tnr_4')
// (15, 24, 'neigh_op_rgt_4')
// (15, 24, 'sp12_h_r_15')
// (15, 25, 'neigh_op_bnr_4')
// (16, 23, 'neigh_op_top_4')
// (16, 24, 'lutff_4/out')
// (16, 24, 'sp12_h_r_16')
// (16, 25, 'neigh_op_bot_4')
// (17, 23, 'neigh_op_tnl_4')
// (17, 24, 'neigh_op_lft_4')
// (17, 24, 'sp12_h_r_19')
// (17, 25, 'neigh_op_bnl_4')
// (18, 24, 'sp12_h_r_20')
// (19, 24, 'sp12_h_r_23')
// (20, 24, 'sp12_h_l_23')
// (20, 24, 'sp12_h_r_0')
// (21, 24, 'sp12_h_r_3')
// (22, 24, 'sp12_h_r_4')
// (23, 24, 'sp12_h_r_7')
// (24, 24, 'sp12_h_r_8')
// (25, 24, 'sp12_h_r_11')
// (26, 24, 'sp12_h_r_12')
// (27, 24, 'sp12_h_r_15')
// (28, 24, 'sp12_h_r_16')
// (29, 24, 'sp12_h_r_19')
// (30, 24, 'sp12_h_r_20')
// (31, 7, 'sp4_r_v_b_47')
// (31, 8, 'sp4_r_v_b_34')
// (31, 9, 'sp4_r_v_b_23')
// (31, 10, 'sp4_r_v_b_10')
// (31, 11, 'sp4_r_v_b_47')
// (31, 12, 'sp4_r_v_b_34')
// (31, 13, 'sp4_r_v_b_23')
// (31, 14, 'sp4_r_v_b_10')
// (31, 24, 'sp12_h_r_23')
// (32, 6, 'sp4_h_r_3')
// (32, 6, 'sp4_v_t_47')
// (32, 7, 'sp4_v_b_47')
// (32, 8, 'sp4_v_b_34')
// (32, 9, 'sp4_v_b_23')
// (32, 10, 'sp4_v_b_10')
// (32, 10, 'sp4_v_t_47')
// (32, 11, 'sp4_v_b_47')
// (32, 12, 'sp12_v_t_23')
// (32, 12, 'sp4_v_b_34')
// (32, 13, 'sp12_v_b_23')
// (32, 13, 'sp4_v_b_23')
// (32, 14, 'sp12_v_b_20')
// (32, 14, 'sp4_v_b_10')
// (32, 15, 'sp12_v_b_19')
// (32, 16, 'sp12_v_b_16')
// (32, 17, 'sp12_v_b_15')
// (32, 18, 'sp12_v_b_12')
// (32, 19, 'sp12_v_b_11')
// (32, 20, 'sp12_v_b_8')
// (32, 21, 'sp12_v_b_7')
// (32, 22, 'sp12_v_b_4')
// (32, 23, 'sp12_v_b_3')
// (32, 24, 'sp12_h_l_23')
// (32, 24, 'sp12_v_b_0')
// (33, 6, 'io_1/D_OUT_0')
// (33, 6, 'local_g0_3')
// (33, 6, 'span4_horz_3')

reg io_11_33_1 = 0;
// (8, 28, 'sp12_h_r_0')
// (9, 28, 'sp12_h_r_3')
// (10, 28, 'sp12_h_r_4')
// (10, 29, 'sp4_r_v_b_40')
// (10, 30, 'sp4_r_v_b_29')
// (10, 31, 'sp4_r_v_b_16')
// (10, 32, 'sp4_r_v_b_5')
// (11, 28, 'sp12_h_r_7')
// (11, 28, 'sp4_h_r_5')
// (11, 28, 'sp4_v_t_40')
// (11, 29, 'sp4_v_b_40')
// (11, 30, 'sp4_v_b_29')
// (11, 31, 'sp4_v_b_16')
// (11, 32, 'sp4_v_b_5')
// (11, 32, 'sp4_v_t_45')
// (11, 33, 'io_1/D_OUT_0')
// (11, 33, 'io_1/PAD')
// (11, 33, 'local_g0_5')
// (11, 33, 'span4_vert_45')
// (12, 28, 'sp12_h_r_8')
// (12, 28, 'sp4_h_r_16')
// (13, 28, 'sp12_h_r_11')
// (13, 28, 'sp4_h_r_29')
// (14, 28, 'sp12_h_r_12')
// (14, 28, 'sp4_h_r_40')
// (15, 28, 'sp12_h_r_15')
// (15, 28, 'sp4_h_l_40')
// (16, 20, 'local_g0_2')
// (16, 20, 'lutff_0/in_2')
// (16, 20, 'sp4_h_r_10')
// (16, 28, 'sp12_h_r_16')
// (17, 20, 'sp4_h_r_23')
// (17, 28, 'sp12_h_r_19')
// (18, 20, 'sp4_h_r_34')
// (18, 22, 'sp12_h_r_0')
// (18, 28, 'sp12_h_r_20')
// (19, 20, 'sp4_h_r_47')
// (19, 21, 'neigh_op_tnr_6')
// (19, 21, 'sp4_r_v_b_41')
// (19, 22, 'neigh_op_rgt_6')
// (19, 22, 'sp12_h_r_3')
// (19, 22, 'sp4_r_v_b_28')
// (19, 23, 'neigh_op_bnr_6')
// (19, 23, 'sp4_r_v_b_17')
// (19, 24, 'sp4_r_v_b_4')
// (19, 28, 'sp12_h_r_23')
// (20, 16, 'sp12_v_t_23')
// (20, 17, 'sp12_v_b_23')
// (20, 18, 'sp12_v_b_20')
// (20, 19, 'sp12_v_b_19')
// (20, 20, 'sp12_v_b_16')
// (20, 20, 'sp4_h_l_47')
// (20, 20, 'sp4_v_t_41')
// (20, 21, 'neigh_op_top_6')
// (20, 21, 'sp12_v_b_15')
// (20, 21, 'sp4_v_b_41')
// (20, 22, 'local_g2_6')
// (20, 22, 'lutff_6/in_0')
// (20, 22, 'lutff_6/out')
// (20, 22, 'lutff_7/in_3')
// (20, 22, 'sp12_h_r_4')
// (20, 22, 'sp12_v_b_12')
// (20, 22, 'sp4_v_b_28')
// (20, 23, 'neigh_op_bot_6')
// (20, 23, 'sp12_v_b_11')
// (20, 23, 'sp4_v_b_17')
// (20, 24, 'sp12_v_b_8')
// (20, 24, 'sp4_v_b_4')
// (20, 25, 'sp12_v_b_7')
// (20, 26, 'sp12_v_b_4')
// (20, 27, 'sp12_v_b_3')
// (20, 28, 'sp12_h_l_23')
// (20, 28, 'sp12_v_b_0')
// (21, 21, 'neigh_op_tnl_6')
// (21, 22, 'neigh_op_lft_6')
// (21, 22, 'sp12_h_r_7')
// (21, 23, 'neigh_op_bnl_6')
// (22, 22, 'sp12_h_r_8')
// (23, 22, 'sp12_h_r_11')
// (24, 22, 'local_g0_4')
// (24, 22, 'lutff_4/in_0')
// (24, 22, 'sp12_h_r_12')
// (25, 22, 'sp12_h_r_15')
// (26, 22, 'sp12_h_r_16')
// (27, 22, 'sp12_h_r_19')
// (28, 22, 'sp12_h_r_20')
// (29, 22, 'sp12_h_r_23')
// (30, 22, 'sp12_h_l_23')

reg n194 = 0;
// (9, 8, 'neigh_op_tnr_0')
// (9, 9, 'neigh_op_rgt_0')
// (9, 10, 'neigh_op_bnr_0')
// (10, 8, 'neigh_op_top_0')
// (10, 9, 'local_g3_0')
// (10, 9, 'lutff_0/in_1')
// (10, 9, 'lutff_0/out')
// (10, 10, 'local_g0_0')
// (10, 10, 'lutff_0/in_2')
// (10, 10, 'neigh_op_bot_0')
// (11, 8, 'neigh_op_tnl_0')
// (11, 9, 'local_g0_0')
// (11, 9, 'lutff_3/in_1')
// (11, 9, 'neigh_op_lft_0')
// (11, 10, 'local_g3_0')
// (11, 10, 'lutff_5/in_2')
// (11, 10, 'neigh_op_bnl_0')

reg n195 = 0;
// (9, 8, 'neigh_op_tnr_1')
// (9, 9, 'neigh_op_rgt_1')
// (9, 9, 'sp4_h_r_7')
// (9, 10, 'neigh_op_bnr_1')
// (10, 8, 'neigh_op_top_1')
// (10, 9, 'local_g0_1')
// (10, 9, 'lutff_1/in_2')
// (10, 9, 'lutff_1/out')
// (10, 9, 'sp4_h_r_18')
// (10, 10, 'local_g1_1')
// (10, 10, 'lutff_1/in_1')
// (10, 10, 'neigh_op_bot_1')
// (11, 8, 'neigh_op_tnl_1')
// (11, 9, 'local_g1_1')
// (11, 9, 'lutff_3/in_3')
// (11, 9, 'neigh_op_lft_1')
// (11, 9, 'sp4_h_r_31')
// (11, 10, 'neigh_op_bnl_1')
// (12, 9, 'sp4_h_r_42')
// (12, 10, 'local_g3_2')
// (12, 10, 'lutff_3/in_0')
// (12, 10, 'sp4_r_v_b_42')
// (12, 11, 'sp4_r_v_b_31')
// (12, 12, 'sp4_r_v_b_18')
// (12, 13, 'sp4_r_v_b_7')
// (13, 9, 'sp4_h_l_42')
// (13, 9, 'sp4_h_r_7')
// (13, 9, 'sp4_v_t_42')
// (13, 10, 'sp4_v_b_42')
// (13, 11, 'sp4_v_b_31')
// (13, 12, 'sp4_v_b_18')
// (13, 13, 'sp4_v_b_7')
// (14, 9, 'local_g1_2')
// (14, 9, 'lutff_5/in_0')
// (14, 9, 'sp4_h_r_18')
// (15, 9, 'sp4_h_r_31')
// (16, 9, 'sp4_h_r_42')
// (17, 9, 'sp4_h_l_42')

reg n196 = 0;
// (9, 8, 'neigh_op_tnr_3')
// (9, 9, 'neigh_op_rgt_3')
// (9, 9, 'sp4_r_v_b_38')
// (9, 10, 'neigh_op_bnr_3')
// (9, 10, 'sp4_r_v_b_27')
// (9, 11, 'sp4_r_v_b_14')
// (9, 12, 'sp4_r_v_b_3')
// (10, 8, 'neigh_op_top_3')
// (10, 8, 'sp4_v_t_38')
// (10, 9, 'lutff_3/out')
// (10, 9, 'sp4_v_b_38')
// (10, 10, 'neigh_op_bot_3')
// (10, 10, 'sp4_v_b_27')
// (10, 11, 'sp4_v_b_14')
// (10, 12, 'local_g0_3')
// (10, 12, 'lutff_1/in_0')
// (10, 12, 'sp4_v_b_3')
// (11, 8, 'neigh_op_tnl_3')
// (11, 9, 'neigh_op_lft_3')
// (11, 10, 'neigh_op_bnl_3')

wire n197;
// (9, 9, 'neigh_op_tnr_1')
// (9, 10, 'neigh_op_rgt_1')
// (9, 11, 'neigh_op_bnr_1')
// (10, 9, 'local_g1_1')
// (10, 9, 'lutff_1/in_1')
// (10, 9, 'neigh_op_top_1')
// (10, 10, 'lutff_1/out')
// (10, 11, 'neigh_op_bot_1')
// (11, 9, 'neigh_op_tnl_1')
// (11, 10, 'neigh_op_lft_1')
// (11, 11, 'neigh_op_bnl_1')

wire n198;
// (9, 9, 'neigh_op_tnr_2')
// (9, 10, 'neigh_op_rgt_2')
// (9, 11, 'neigh_op_bnr_2')
// (10, 9, 'neigh_op_top_2')
// (10, 10, 'lutff_2/out')
// (10, 11, 'neigh_op_bot_2')
// (11, 9, 'local_g2_2')
// (11, 9, 'lutff_7/in_3')
// (11, 9, 'neigh_op_tnl_2')
// (11, 10, 'neigh_op_lft_2')
// (11, 11, 'neigh_op_bnl_2')

wire n199;
// (9, 9, 'neigh_op_tnr_3')
// (9, 10, 'neigh_op_rgt_3')
// (9, 11, 'neigh_op_bnr_3')
// (10, 9, 'local_g1_3')
// (10, 9, 'lutff_5/in_3')
// (10, 9, 'neigh_op_top_3')
// (10, 10, 'lutff_3/out')
// (10, 11, 'neigh_op_bot_3')
// (11, 9, 'neigh_op_tnl_3')
// (11, 10, 'neigh_op_lft_3')
// (11, 11, 'neigh_op_bnl_3')

reg n200 = 0;
// (9, 9, 'neigh_op_tnr_4')
// (9, 10, 'neigh_op_rgt_4')
// (9, 11, 'neigh_op_bnr_4')
// (10, 9, 'neigh_op_top_4')
// (10, 10, 'local_g3_4')
// (10, 10, 'lutff_4/in_1')
// (10, 10, 'lutff_4/out')
// (10, 11, 'neigh_op_bot_4')
// (11, 9, 'local_g3_4')
// (11, 9, 'lutff_3/in_0')
// (11, 9, 'neigh_op_tnl_4')
// (11, 10, 'neigh_op_lft_4')
// (11, 11, 'neigh_op_bnl_4')

reg n201 = 0;
// (9, 10, 'neigh_op_tnr_0')
// (9, 11, 'neigh_op_rgt_0')
// (9, 12, 'neigh_op_bnr_0')
// (10, 9, 'sp4_r_v_b_41')
// (10, 10, 'neigh_op_top_0')
// (10, 10, 'sp4_r_v_b_28')
// (10, 11, 'local_g1_0')
// (10, 11, 'lutff_0/in_1')
// (10, 11, 'lutff_0/out')
// (10, 11, 'sp4_r_v_b_17')
// (10, 12, 'neigh_op_bot_0')
// (10, 12, 'sp4_r_v_b_4')
// (11, 8, 'sp4_v_t_41')
// (11, 9, 'local_g2_1')
// (11, 9, 'lutff_3/in_2')
// (11, 9, 'sp4_v_b_41')
// (11, 10, 'neigh_op_tnl_0')
// (11, 10, 'sp4_v_b_28')
// (11, 11, 'neigh_op_lft_0')
// (11, 11, 'sp4_v_b_17')
// (11, 12, 'neigh_op_bnl_0')
// (11, 12, 'sp4_v_b_4')

reg n202 = 0;
// (9, 11, 'sp12_h_r_1')
// (10, 11, 'sp12_h_r_2')
// (11, 11, 'sp12_h_r_5')
// (12, 11, 'sp12_h_r_6')
// (13, 11, 'sp12_h_r_9')
// (14, 11, 'sp12_h_r_10')
// (15, 10, 'neigh_op_tnr_3')
// (15, 11, 'neigh_op_rgt_3')
// (15, 11, 'sp12_h_r_13')
// (15, 12, 'neigh_op_bnr_3')
// (16, 10, 'neigh_op_top_3')
// (16, 11, 'lutff_3/out')
// (16, 11, 'sp12_h_r_14')
// (16, 12, 'neigh_op_bot_3')
// (17, 10, 'neigh_op_tnl_3')
// (17, 11, 'neigh_op_lft_3')
// (17, 11, 'sp12_h_r_17')
// (17, 12, 'neigh_op_bnl_3')
// (18, 11, 'sp12_h_r_18')
// (19, 11, 'sp12_h_r_21')
// (20, 11, 'sp12_h_r_22')
// (21, 11, 'sp12_h_l_22')
// (21, 11, 'sp12_v_t_22')
// (21, 12, 'sp12_v_b_22')
// (21, 13, 'sp12_v_b_21')
// (21, 14, 'sp12_v_b_18')
// (21, 15, 'local_g2_1')
// (21, 15, 'lutff_0/in_1')
// (21, 15, 'sp12_v_b_17')
// (21, 16, 'sp12_v_b_14')
// (21, 17, 'sp12_v_b_13')
// (21, 18, 'sp12_v_b_10')
// (21, 19, 'sp12_v_b_9')
// (21, 20, 'sp12_v_b_6')
// (21, 21, 'sp12_v_b_5')
// (21, 22, 'sp12_v_b_2')
// (21, 23, 'sp12_v_b_1')

reg n203 = 0;
// (9, 12, 'local_g2_0')
// (9, 12, 'lutff_5/in_3')
// (9, 12, 'neigh_op_tnr_0')
// (9, 13, 'neigh_op_rgt_0')
// (9, 14, 'neigh_op_bnr_0')
// (10, 12, 'neigh_op_top_0')
// (10, 13, 'local_g3_0')
// (10, 13, 'lutff_0/in_1')
// (10, 13, 'lutff_0/out')
// (10, 14, 'neigh_op_bot_0')
// (11, 12, 'neigh_op_tnl_0')
// (11, 13, 'neigh_op_lft_0')
// (11, 14, 'neigh_op_bnl_0')

reg n204 = 0;
// (9, 12, 'local_g3_4')
// (9, 12, 'lutff_5/in_0')
// (9, 12, 'neigh_op_tnr_4')
// (9, 13, 'neigh_op_rgt_4')
// (9, 14, 'neigh_op_bnr_4')
// (10, 12, 'neigh_op_top_4')
// (10, 13, 'local_g3_4')
// (10, 13, 'lutff_4/in_1')
// (10, 13, 'lutff_4/out')
// (10, 14, 'neigh_op_bot_4')
// (11, 12, 'neigh_op_tnl_4')
// (11, 13, 'neigh_op_lft_4')
// (11, 14, 'neigh_op_bnl_4')

wire n205;
// (9, 12, 'lutff_2/lout')
// (9, 12, 'lutff_3/in_2')

reg n206 = 0;
// (9, 12, 'neigh_op_tnr_1')
// (9, 13, 'neigh_op_rgt_1')
// (9, 14, 'local_g0_1')
// (9, 14, 'lutff_7/in_0')
// (9, 14, 'neigh_op_bnr_1')
// (10, 12, 'neigh_op_top_1')
// (10, 13, 'local_g3_1')
// (10, 13, 'lutff_1/in_1')
// (10, 13, 'lutff_1/out')
// (10, 14, 'neigh_op_bot_1')
// (11, 12, 'neigh_op_tnl_1')
// (11, 13, 'neigh_op_lft_1')
// (11, 14, 'neigh_op_bnl_1')

reg n207 = 0;
// (9, 12, 'neigh_op_tnr_2')
// (9, 13, 'neigh_op_rgt_2')
// (9, 14, 'local_g1_2')
// (9, 14, 'lutff_7/in_2')
// (9, 14, 'neigh_op_bnr_2')
// (10, 12, 'neigh_op_top_2')
// (10, 13, 'local_g1_2')
// (10, 13, 'lutff_2/in_1')
// (10, 13, 'lutff_2/out')
// (10, 14, 'neigh_op_bot_2')
// (11, 12, 'neigh_op_tnl_2')
// (11, 13, 'neigh_op_lft_2')
// (11, 14, 'neigh_op_bnl_2')

reg n208 = 0;
// (9, 12, 'neigh_op_tnr_3')
// (9, 13, 'neigh_op_rgt_3')
// (9, 14, 'neigh_op_bnr_3')
// (10, 12, 'neigh_op_top_3')
// (10, 13, 'local_g1_3')
// (10, 13, 'lutff_3/in_1')
// (10, 13, 'lutff_3/out')
// (10, 14, 'local_g1_3')
// (10, 14, 'lutff_7/in_3')
// (10, 14, 'neigh_op_bot_3')
// (11, 12, 'neigh_op_tnl_3')
// (11, 13, 'neigh_op_lft_3')
// (11, 14, 'neigh_op_bnl_3')

reg n209 = 0;
// (9, 12, 'neigh_op_tnr_5')
// (9, 13, 'neigh_op_rgt_5')
// (9, 14, 'neigh_op_bnr_5')
// (10, 12, 'neigh_op_top_5')
// (10, 13, 'local_g1_5')
// (10, 13, 'lutff_5/in_1')
// (10, 13, 'lutff_5/out')
// (10, 14, 'local_g1_5')
// (10, 14, 'lutff_7/in_1')
// (10, 14, 'neigh_op_bot_5')
// (11, 12, 'neigh_op_tnl_5')
// (11, 13, 'neigh_op_lft_5')
// (11, 14, 'neigh_op_bnl_5')

reg n210 = 0;
// (9, 12, 'neigh_op_tnr_6')
// (9, 13, 'neigh_op_rgt_6')
// (9, 14, 'neigh_op_bnr_6')
// (10, 12, 'neigh_op_top_6')
// (10, 13, 'local_g1_6')
// (10, 13, 'lutff_6/in_1')
// (10, 13, 'lutff_6/out')
// (10, 14, 'local_g1_6')
// (10, 14, 'lutff_7/in_0')
// (10, 14, 'neigh_op_bot_6')
// (11, 12, 'neigh_op_tnl_6')
// (11, 13, 'neigh_op_lft_6')
// (11, 14, 'neigh_op_bnl_6')

reg n211 = 0;
// (9, 12, 'neigh_op_tnr_7')
// (9, 13, 'neigh_op_rgt_7')
// (9, 14, 'neigh_op_bnr_7')
// (10, 12, 'neigh_op_top_7')
// (10, 13, 'local_g2_7')
// (10, 13, 'lutff_7/in_0')
// (10, 13, 'lutff_7/out')
// (10, 14, 'local_g0_7')
// (10, 14, 'lutff_7/in_2')
// (10, 14, 'neigh_op_bot_7')
// (11, 12, 'neigh_op_tnl_7')
// (11, 13, 'neigh_op_lft_7')
// (11, 14, 'neigh_op_bnl_7')

reg n212 = 0;
// (9, 12, 'sp4_h_r_10')
// (9, 13, 'sp4_r_v_b_36')
// (9, 14, 'sp4_r_v_b_25')
// (9, 15, 'sp4_r_v_b_12')
// (9, 16, 'local_g1_1')
// (9, 16, 'lutff_7/in_3')
// (9, 16, 'sp4_r_v_b_1')
// (9, 17, 'local_g3_1')
// (9, 17, 'lutff_5/in_3')
// (9, 17, 'sp4_r_v_b_41')
// (9, 18, 'sp4_r_v_b_28')
// (9, 19, 'sp4_r_v_b_17')
// (9, 20, 'sp4_r_v_b_4')
// (10, 11, 'neigh_op_tnr_1')
// (10, 12, 'neigh_op_rgt_1')
// (10, 12, 'sp4_h_r_23')
// (10, 12, 'sp4_h_r_7')
// (10, 12, 'sp4_v_t_36')
// (10, 13, 'neigh_op_bnr_1')
// (10, 13, 'sp4_v_b_36')
// (10, 14, 'sp4_v_b_25')
// (10, 15, 'sp4_v_b_12')
// (10, 16, 'sp4_v_b_1')
// (10, 16, 'sp4_v_t_41')
// (10, 17, 'sp4_v_b_41')
// (10, 18, 'sp4_v_b_28')
// (10, 19, 'local_g1_1')
// (10, 19, 'lutff_1/in_3')
// (10, 19, 'sp4_v_b_17')
// (10, 20, 'local_g0_4')
// (10, 20, 'lutff_7/in_3')
// (10, 20, 'sp4_v_b_4')
// (11, 9, 'sp12_v_t_22')
// (11, 10, 'sp12_v_b_22')
// (11, 11, 'neigh_op_top_1')
// (11, 11, 'sp12_v_b_21')
// (11, 12, 'lutff_1/out')
// (11, 12, 'sp12_v_b_18')
// (11, 12, 'sp4_h_r_18')
// (11, 12, 'sp4_h_r_2')
// (11, 12, 'sp4_h_r_34')
// (11, 13, 'local_g1_1')
// (11, 13, 'lutff_7/in_3')
// (11, 13, 'neigh_op_bot_1')
// (11, 13, 'sp12_v_b_17')
// (11, 14, 'sp12_v_b_14')
// (11, 15, 'sp12_v_b_13')
// (11, 16, 'sp12_v_b_10')
// (11, 17, 'sp12_v_b_9')
// (11, 18, 'sp12_v_b_6')
// (11, 19, 'sp12_v_b_5')
// (11, 20, 'sp12_v_b_2')
// (11, 21, 'sp12_h_r_1')
// (11, 21, 'sp12_v_b_1')
// (11, 21, 'sp12_v_t_22')
// (11, 22, 'local_g2_6')
// (11, 22, 'lutff_1/in_3')
// (11, 22, 'sp12_v_b_22')
// (11, 23, 'sp12_v_b_21')
// (11, 24, 'sp12_v_b_18')
// (11, 25, 'sp12_v_b_17')
// (11, 26, 'sp12_v_b_14')
// (11, 27, 'sp12_v_b_13')
// (11, 28, 'sp12_v_b_10')
// (11, 29, 'sp12_v_b_9')
// (11, 30, 'sp12_v_b_6')
// (11, 31, 'sp12_v_b_5')
// (11, 32, 'sp12_v_b_2')
// (11, 33, 'span12_vert_1')
// (12, 11, 'neigh_op_tnl_1')
// (12, 12, 'neigh_op_lft_1')
// (12, 12, 'sp4_h_r_15')
// (12, 12, 'sp4_h_r_31')
// (12, 12, 'sp4_h_r_47')
// (12, 13, 'local_g3_1')
// (12, 13, 'lutff_1/in_3')
// (12, 13, 'neigh_op_bnl_1')
// (12, 13, 'sp4_r_v_b_38')
// (12, 14, 'sp4_r_v_b_27')
// (12, 15, 'sp4_r_v_b_14')
// (12, 16, 'sp4_r_v_b_3')
// (12, 17, 'sp4_r_v_b_38')
// (12, 18, 'sp4_r_v_b_27')
// (12, 19, 'local_g2_6')
// (12, 19, 'lutff_1/in_3')
// (12, 19, 'sp4_r_v_b_14')
// (12, 20, 'sp4_r_v_b_3')
// (12, 21, 'sp12_h_r_2')
// (13, 12, 'sp4_h_l_47')
// (13, 12, 'sp4_h_r_1')
// (13, 12, 'sp4_h_r_26')
// (13, 12, 'sp4_h_r_42')
// (13, 12, 'sp4_v_t_38')
// (13, 13, 'sp4_r_v_b_37')
// (13, 13, 'sp4_v_b_38')
// (13, 14, 'sp4_r_v_b_24')
// (13, 14, 'sp4_v_b_27')
// (13, 15, 'sp4_r_v_b_13')
// (13, 15, 'sp4_v_b_14')
// (13, 16, 'local_g1_0')
// (13, 16, 'lutff_7/in_0')
// (13, 16, 'sp4_h_r_3')
// (13, 16, 'sp4_r_v_b_0')
// (13, 16, 'sp4_v_b_3')
// (13, 16, 'sp4_v_t_38')
// (13, 17, 'sp4_v_b_38')
// (13, 18, 'sp4_v_b_27')
// (13, 19, 'sp4_v_b_14')
// (13, 20, 'sp4_v_b_3')
// (13, 21, 'sp12_h_r_5')
// (14, 12, 'sp4_h_l_42')
// (14, 12, 'sp4_h_r_10')
// (14, 12, 'sp4_h_r_12')
// (14, 12, 'sp4_h_r_39')
// (14, 12, 'sp4_v_t_37')
// (14, 13, 'local_g3_5')
// (14, 13, 'lutff_1/in_3')
// (14, 13, 'sp4_r_v_b_39')
// (14, 13, 'sp4_v_b_37')
// (14, 14, 'sp4_r_v_b_26')
// (14, 14, 'sp4_v_b_24')
// (14, 15, 'sp4_r_v_b_15')
// (14, 15, 'sp4_v_b_13')
// (14, 16, 'sp4_h_r_14')
// (14, 16, 'sp4_r_v_b_2')
// (14, 16, 'sp4_v_b_0')
// (14, 17, 'sp4_r_v_b_47')
// (14, 18, 'sp4_r_v_b_34')
// (14, 19, 'sp4_r_v_b_23')
// (14, 20, 'sp4_r_v_b_10')
// (14, 21, 'sp12_h_r_6')
// (14, 21, 'sp4_r_v_b_36')
// (14, 22, 'sp4_r_v_b_25')
// (14, 23, 'local_g2_4')
// (14, 23, 'lutff_7/in_3')
// (14, 23, 'sp4_r_v_b_12')
// (14, 24, 'sp4_r_v_b_1')
// (15, 12, 'sp4_h_l_39')
// (15, 12, 'sp4_h_r_23')
// (15, 12, 'sp4_h_r_25')
// (15, 12, 'sp4_h_r_5')
// (15, 12, 'sp4_v_t_39')
// (15, 13, 'sp4_v_b_39')
// (15, 14, 'sp4_v_b_26')
// (15, 15, 'local_g1_7')
// (15, 15, 'lutff_1/in_3')
// (15, 15, 'sp4_v_b_15')
// (15, 16, 'sp4_h_r_27')
// (15, 16, 'sp4_v_b_2')
// (15, 16, 'sp4_v_t_47')
// (15, 17, 'local_g3_7')
// (15, 17, 'lutff_1/in_3')
// (15, 17, 'sp4_v_b_47')
// (15, 18, 'local_g3_2')
// (15, 18, 'lutff_1/in_0')
// (15, 18, 'sp4_v_b_34')
// (15, 19, 'local_g1_7')
// (15, 19, 'lutff_1/in_3')
// (15, 19, 'sp4_v_b_23')
// (15, 20, 'sp4_v_b_10')
// (15, 20, 'sp4_v_t_36')
// (15, 21, 'sp12_h_r_9')
// (15, 21, 'sp4_h_r_4')
// (15, 21, 'sp4_v_b_36')
// (15, 22, 'sp4_v_b_25')
// (15, 23, 'sp4_v_b_12')
// (15, 24, 'sp4_v_b_1')
// (16, 9, 'sp4_r_v_b_36')
// (16, 10, 'sp4_r_v_b_25')
// (16, 11, 'local_g2_4')
// (16, 11, 'lutff_1/in_3')
// (16, 11, 'sp4_r_v_b_12')
// (16, 12, 'local_g2_2')
// (16, 12, 'lutff_1/in_1')
// (16, 12, 'sp4_h_r_16')
// (16, 12, 'sp4_h_r_34')
// (16, 12, 'sp4_h_r_36')
// (16, 12, 'sp4_r_v_b_1')
// (16, 16, 'local_g2_6')
// (16, 16, 'lutff_1/in_3')
// (16, 16, 'sp4_h_r_38')
// (16, 17, 'local_g2_6')
// (16, 17, 'lutff_1/in_3')
// (16, 17, 'sp4_r_v_b_38')
// (16, 18, 'local_g0_3')
// (16, 18, 'lutff_1/in_0')
// (16, 18, 'sp4_r_v_b_27')
// (16, 19, 'local_g2_6')
// (16, 19, 'lutff_7/in_3')
// (16, 19, 'sp4_r_v_b_14')
// (16, 20, 'sp4_r_v_b_3')
// (16, 21, 'local_g0_2')
// (16, 21, 'lutff_7/in_3')
// (16, 21, 'sp12_h_r_10')
// (16, 21, 'sp4_h_r_17')
// (17, 8, 'sp4_v_t_36')
// (17, 9, 'sp4_r_v_b_41')
// (17, 9, 'sp4_v_b_36')
// (17, 10, 'sp4_r_v_b_28')
// (17, 10, 'sp4_v_b_25')
// (17, 11, 'sp4_r_v_b_17')
// (17, 11, 'sp4_v_b_12')
// (17, 12, 'sp4_h_l_36')
// (17, 12, 'sp4_h_r_29')
// (17, 12, 'sp4_h_r_47')
// (17, 12, 'sp4_h_r_9')
// (17, 12, 'sp4_r_v_b_4')
// (17, 12, 'sp4_v_b_1')
// (17, 16, 'sp4_h_l_38')
// (17, 16, 'sp4_v_t_38')
// (17, 17, 'local_g3_6')
// (17, 17, 'lutff_4/in_3')
// (17, 17, 'sp4_v_b_38')
// (17, 18, 'sp4_v_b_27')
// (17, 19, 'sp4_v_b_14')
// (17, 20, 'sp4_v_b_3')
// (17, 21, 'sp12_h_r_13')
// (17, 21, 'sp4_h_r_28')
// (18, 8, 'sp4_v_t_41')
// (18, 9, 'sp4_r_v_b_46')
// (18, 9, 'sp4_v_b_41')
// (18, 10, 'sp4_r_v_b_35')
// (18, 10, 'sp4_v_b_28')
// (18, 11, 'local_g1_1')
// (18, 11, 'lutff_1/in_3')
// (18, 11, 'sp4_r_v_b_22')
// (18, 11, 'sp4_v_b_17')
// (18, 12, 'local_g0_4')
// (18, 12, 'lutff_1/in_3')
// (18, 12, 'sp4_h_l_47')
// (18, 12, 'sp4_h_r_1')
// (18, 12, 'sp4_h_r_20')
// (18, 12, 'sp4_h_r_40')
// (18, 12, 'sp4_r_v_b_11')
// (18, 12, 'sp4_v_b_4')
// (18, 13, 'sp4_r_v_b_47')
// (18, 14, 'sp4_r_v_b_34')
// (18, 15, 'sp4_r_v_b_23')
// (18, 16, 'sp4_r_v_b_10')
// (18, 21, 'sp12_h_r_14')
// (18, 21, 'sp4_h_r_41')
// (18, 22, 'sp4_r_v_b_41')
// (18, 23, 'sp4_r_v_b_28')
// (18, 24, 'sp4_r_v_b_17')
// (18, 25, 'sp4_r_v_b_4')
// (19, 8, 'sp4_v_t_46')
// (19, 9, 'sp4_v_b_46')
// (19, 10, 'local_g3_3')
// (19, 10, 'lutff_1/in_3')
// (19, 10, 'sp4_v_b_35')
// (19, 11, 'local_g0_6')
// (19, 11, 'lutff_1/in_3')
// (19, 11, 'sp4_v_b_22')
// (19, 12, 'sp4_h_l_40')
// (19, 12, 'sp4_h_r_12')
// (19, 12, 'sp4_h_r_33')
// (19, 12, 'sp4_h_r_5')
// (19, 12, 'sp4_v_b_11')
// (19, 12, 'sp4_v_t_47')
// (19, 13, 'sp4_v_b_47')
// (19, 14, 'sp4_v_b_34')
// (19, 15, 'local_g0_7')
// (19, 15, 'lutff_5/in_0')
// (19, 15, 'sp4_v_b_23')
// (19, 16, 'local_g0_2')
// (19, 16, 'lutff_1/in_3')
// (19, 16, 'sp4_v_b_10')
// (19, 21, 'sp12_h_r_17')
// (19, 21, 'sp4_h_l_41')
// (19, 21, 'sp4_h_r_8')
// (19, 21, 'sp4_v_t_41')
// (19, 22, 'sp4_v_b_41')
// (19, 23, 'sp4_v_b_28')
// (19, 24, 'sp4_v_b_17')
// (19, 25, 'local_g0_4')
// (19, 25, 'lutff_1/in_3')
// (19, 25, 'sp4_h_r_4')
// (19, 25, 'sp4_v_b_4')
// (20, 9, 'sp4_r_v_b_44')
// (20, 10, 'sp4_r_v_b_33')
// (20, 11, 'local_g3_4')
// (20, 11, 'lutff_0/in_3')
// (20, 11, 'sp4_r_v_b_20')
// (20, 12, 'local_g2_4')
// (20, 12, 'lutff_1/in_3')
// (20, 12, 'sp4_h_r_16')
// (20, 12, 'sp4_h_r_25')
// (20, 12, 'sp4_h_r_44')
// (20, 12, 'sp4_r_v_b_9')
// (20, 13, 'local_g2_7')
// (20, 13, 'lutff_5/in_0')
// (20, 13, 'sp4_r_v_b_39')
// (20, 14, 'sp4_r_v_b_26')
// (20, 15, 'sp4_r_v_b_15')
// (20, 16, 'local_g1_2')
// (20, 16, 'lutff_1/in_0')
// (20, 16, 'sp4_r_v_b_2')
// (20, 17, 'local_g3_0')
// (20, 17, 'lutff_3/in_0')
// (20, 17, 'sp4_r_v_b_40')
// (20, 18, 'local_g0_5')
// (20, 18, 'lutff_4/in_3')
// (20, 18, 'sp4_r_v_b_29')
// (20, 19, 'local_g3_0')
// (20, 19, 'lutff_1/in_0')
// (20, 19, 'sp4_r_v_b_16')
// (20, 20, 'local_g1_5')
// (20, 20, 'lutff_1/in_3')
// (20, 20, 'sp4_r_v_b_5')
// (20, 21, 'sp12_h_r_18')
// (20, 21, 'sp4_h_r_21')
// (20, 21, 'sp4_r_v_b_45')
// (20, 22, 'sp4_r_v_b_32')
// (20, 23, 'local_g3_5')
// (20, 23, 'lutff_3/in_3')
// (20, 23, 'sp4_r_v_b_21')
// (20, 24, 'sp4_r_v_b_8')
// (20, 25, 'local_g1_1')
// (20, 25, 'lutff_1/in_3')
// (20, 25, 'sp4_h_r_17')
// (21, 8, 'sp4_v_t_44')
// (21, 9, 'sp4_v_b_44')
// (21, 10, 'sp4_v_b_33')
// (21, 11, 'local_g0_4')
// (21, 11, 'lutff_1/in_3')
// (21, 11, 'sp4_v_b_20')
// (21, 12, 'local_g2_4')
// (21, 12, 'lutff_1/in_3')
// (21, 12, 'sp4_h_l_44')
// (21, 12, 'sp4_h_r_0')
// (21, 12, 'sp4_h_r_29')
// (21, 12, 'sp4_h_r_36')
// (21, 12, 'sp4_v_b_9')
// (21, 12, 'sp4_v_t_39')
// (21, 13, 'local_g3_7')
// (21, 13, 'lutff_4/in_0')
// (21, 13, 'sp4_r_v_b_43')
// (21, 13, 'sp4_v_b_39')
// (21, 14, 'local_g0_6')
// (21, 14, 'lutff_5/in_3')
// (21, 14, 'sp4_r_v_b_30')
// (21, 14, 'sp4_v_b_26')
// (21, 15, 'sp4_r_v_b_19')
// (21, 15, 'sp4_v_b_15')
// (21, 16, 'sp4_r_v_b_6')
// (21, 16, 'sp4_v_b_2')
// (21, 16, 'sp4_v_t_40')
// (21, 17, 'sp4_v_b_40')
// (21, 18, 'sp4_v_b_29')
// (21, 19, 'sp4_v_b_16')
// (21, 20, 'local_g1_5')
// (21, 20, 'lutff_1/in_3')
// (21, 20, 'sp4_v_b_5')
// (21, 20, 'sp4_v_t_45')
// (21, 21, 'local_g0_5')
// (21, 21, 'lutff_6/in_3')
// (21, 21, 'sp12_h_r_21')
// (21, 21, 'sp4_h_r_32')
// (21, 21, 'sp4_v_b_45')
// (21, 22, 'sp4_v_b_32')
// (21, 23, 'sp4_v_b_21')
// (21, 24, 'sp4_v_b_8')
// (21, 25, 'sp4_h_r_28')
// (22, 12, 'local_g2_0')
// (22, 12, 'lutff_1/in_3')
// (22, 12, 'sp4_h_l_36')
// (22, 12, 'sp4_h_r_13')
// (22, 12, 'sp4_h_r_40')
// (22, 12, 'sp4_v_t_43')
// (22, 13, 'sp4_r_v_b_47')
// (22, 13, 'sp4_v_b_43')
// (22, 14, 'local_g2_6')
// (22, 14, 'lutff_1/in_3')
// (22, 14, 'sp4_r_v_b_34')
// (22, 14, 'sp4_v_b_30')
// (22, 15, 'sp4_r_v_b_23')
// (22, 15, 'sp4_v_b_19')
// (22, 16, 'sp4_r_v_b_10')
// (22, 16, 'sp4_v_b_6')
// (22, 21, 'local_g0_6')
// (22, 21, 'lutff_1/in_3')
// (22, 21, 'sp12_h_r_22')
// (22, 21, 'sp4_h_r_45')
// (22, 22, 'sp4_r_v_b_45')
// (22, 23, 'local_g2_0')
// (22, 23, 'lutff_1/in_3')
// (22, 23, 'sp4_r_v_b_32')
// (22, 24, 'sp4_r_v_b_21')
// (22, 25, 'sp4_h_r_41')
// (22, 25, 'sp4_r_v_b_8')
// (23, 9, 'sp12_v_t_22')
// (23, 10, 'sp12_v_b_22')
// (23, 11, 'sp12_v_b_21')
// (23, 12, 'local_g2_0')
// (23, 12, 'lutff_1/in_3')
// (23, 12, 'sp12_v_b_18')
// (23, 12, 'sp4_h_l_40')
// (23, 12, 'sp4_h_r_24')
// (23, 12, 'sp4_v_t_47')
// (23, 13, 'sp12_v_b_17')
// (23, 13, 'sp4_v_b_47')
// (23, 14, 'local_g2_2')
// (23, 14, 'lutff_1/in_3')
// (23, 14, 'sp12_v_b_14')
// (23, 14, 'sp4_v_b_34')
// (23, 15, 'local_g1_7')
// (23, 15, 'lutff_1/in_3')
// (23, 15, 'sp12_v_b_13')
// (23, 15, 'sp4_v_b_23')
// (23, 16, 'local_g0_2')
// (23, 16, 'lutff_1/in_3')
// (23, 16, 'sp12_v_b_10')
// (23, 16, 'sp4_v_b_10')
// (23, 17, 'sp12_v_b_9')
// (23, 18, 'local_g2_6')
// (23, 18, 'lutff_1/in_3')
// (23, 18, 'sp12_v_b_6')
// (23, 19, 'sp12_v_b_5')
// (23, 20, 'local_g2_2')
// (23, 20, 'lutff_1/in_3')
// (23, 20, 'sp12_v_b_2')
// (23, 21, 'sp12_h_l_22')
// (23, 21, 'sp12_v_b_1')
// (23, 21, 'sp4_h_l_45')
// (23, 21, 'sp4_v_t_45')
// (23, 22, 'sp4_v_b_45')
// (23, 23, 'sp4_v_b_32')
// (23, 24, 'sp4_v_b_21')
// (23, 25, 'sp4_h_l_41')
// (23, 25, 'sp4_v_b_8')
// (24, 12, 'sp4_h_r_37')
// (24, 13, 'sp4_r_v_b_40')
// (24, 14, 'local_g1_5')
// (24, 14, 'lutff_1/in_3')
// (24, 14, 'sp4_r_v_b_29')
// (24, 15, 'local_g3_0')
// (24, 15, 'lutff_1/in_0')
// (24, 15, 'sp4_r_v_b_16')
// (24, 16, 'sp4_r_v_b_5')
// (24, 17, 'local_g2_4')
// (24, 17, 'lutff_1/in_3')
// (24, 17, 'sp4_r_v_b_36')
// (24, 18, 'sp4_r_v_b_25')
// (24, 19, 'sp4_r_v_b_12')
// (24, 20, 'sp4_r_v_b_1')
// (25, 12, 'sp4_h_l_37')
// (25, 12, 'sp4_v_t_40')
// (25, 13, 'sp4_v_b_40')
// (25, 14, 'sp4_v_b_29')
// (25, 15, 'sp4_v_b_16')
// (25, 16, 'sp4_v_b_5')
// (25, 16, 'sp4_v_t_36')
// (25, 17, 'sp4_v_b_36')
// (25, 18, 'sp4_v_b_25')
// (25, 19, 'sp4_v_b_12')
// (25, 20, 'sp4_v_b_1')

reg n213 = 0;
// (9, 13, 'neigh_op_tnr_1')
// (9, 14, 'neigh_op_rgt_1')
// (9, 15, 'local_g1_1')
// (9, 15, 'lutff_1/in_1')
// (9, 15, 'neigh_op_bnr_1')
// (10, 13, 'neigh_op_top_1')
// (10, 14, 'local_g3_1')
// (10, 14, 'lutff_1/in_3')
// (10, 14, 'lutff_1/out')
// (10, 14, 'lutff_2/in_0')
// (10, 15, 'local_g0_1')
// (10, 15, 'lutff_0/in_1')
// (10, 15, 'neigh_op_bot_1')
// (11, 13, 'neigh_op_tnl_1')
// (11, 14, 'neigh_op_lft_1')
// (11, 15, 'neigh_op_bnl_1')

reg n214 = 0;
// (9, 13, 'neigh_op_tnr_2')
// (9, 14, 'neigh_op_rgt_2')
// (9, 15, 'neigh_op_bnr_2')
// (10, 13, 'neigh_op_top_2')
// (10, 14, 'local_g3_2')
// (10, 14, 'lutff_2/in_3')
// (10, 14, 'lutff_2/out')
// (10, 15, 'local_g0_2')
// (10, 15, 'lutff_0/in_2')
// (10, 15, 'neigh_op_bot_2')
// (11, 13, 'neigh_op_tnl_2')
// (11, 14, 'neigh_op_lft_2')
// (11, 15, 'neigh_op_bnl_2')

wire n215;
// (9, 13, 'neigh_op_tnr_3')
// (9, 14, 'neigh_op_rgt_3')
// (9, 15, 'neigh_op_bnr_3')
// (10, 13, 'neigh_op_top_3')
// (10, 14, 'lutff_3/out')
// (10, 14, 'sp4_r_v_b_39')
// (10, 15, 'neigh_op_bot_3')
// (10, 15, 'sp4_r_v_b_26')
// (10, 16, 'sp4_r_v_b_15')
// (10, 17, 'sp4_r_v_b_2')
// (11, 13, 'neigh_op_tnl_3')
// (11, 13, 'sp4_h_r_7')
// (11, 13, 'sp4_v_t_39')
// (11, 14, 'neigh_op_lft_3')
// (11, 14, 'sp4_v_b_39')
// (11, 15, 'neigh_op_bnl_3')
// (11, 15, 'sp4_v_b_26')
// (11, 16, 'sp4_v_b_15')
// (11, 17, 'sp4_v_b_2')
// (12, 13, 'sp4_h_r_18')
// (13, 13, 'sp4_h_r_31')
// (14, 10, 'sp4_r_v_b_42')
// (14, 11, 'sp4_r_v_b_31')
// (14, 12, 'sp4_r_v_b_18')
// (14, 13, 'sp4_h_r_42')
// (14, 13, 'sp4_r_v_b_7')
// (15, 9, 'sp4_h_r_7')
// (15, 9, 'sp4_v_t_42')
// (15, 10, 'sp4_v_b_42')
// (15, 11, 'sp4_v_b_31')
// (15, 12, 'sp4_v_b_18')
// (15, 13, 'sp4_h_l_42')
// (15, 13, 'sp4_v_b_7')
// (16, 9, 'sp4_h_r_18')
// (17, 9, 'sp4_h_r_31')
// (18, 9, 'local_g2_2')
// (18, 9, 'lutff_global/cen')
// (18, 9, 'sp4_h_r_42')
// (19, 9, 'sp4_h_l_42')

wire n216;
// (9, 13, 'neigh_op_tnr_7')
// (9, 14, 'local_g3_7')
// (9, 14, 'lutff_7/in_1')
// (9, 14, 'neigh_op_rgt_7')
// (9, 15, 'neigh_op_bnr_7')
// (10, 13, 'neigh_op_top_7')
// (10, 14, 'lutff_7/out')
// (10, 15, 'neigh_op_bot_7')
// (11, 13, 'neigh_op_tnl_7')
// (11, 14, 'neigh_op_lft_7')
// (11, 15, 'neigh_op_bnl_7')

reg n217 = 0;
// (9, 13, 'sp12_h_r_1')
// (10, 13, 'sp12_h_r_2')
// (11, 13, 'sp12_h_r_5')
// (12, 13, 'sp12_h_r_6')
// (13, 12, 'neigh_op_tnr_1')
// (13, 13, 'neigh_op_rgt_1')
// (13, 13, 'sp12_h_r_9')
// (13, 14, 'neigh_op_bnr_1')
// (14, 12, 'neigh_op_top_1')
// (14, 13, 'lutff_1/out')
// (14, 13, 'sp12_h_r_10')
// (14, 14, 'neigh_op_bot_1')
// (15, 12, 'neigh_op_tnl_1')
// (15, 13, 'neigh_op_lft_1')
// (15, 13, 'sp12_h_r_13')
// (15, 14, 'neigh_op_bnl_1')
// (16, 13, 'sp12_h_r_14')
// (17, 13, 'sp12_h_r_17')
// (18, 13, 'sp12_h_r_18')
// (19, 13, 'local_g0_5')
// (19, 13, 'lutff_4/in_1')
// (19, 13, 'sp12_h_r_21')
// (20, 13, 'sp12_h_r_22')
// (21, 13, 'sp12_h_l_22')

reg n218 = 0;
// (9, 13, 'sp4_r_v_b_44')
// (9, 14, 'sp4_r_v_b_33')
// (9, 15, 'sp4_r_v_b_20')
// (9, 16, 'local_g2_1')
// (9, 16, 'lutff_7/in_2')
// (9, 16, 'sp4_r_v_b_9')
// (9, 17, 'sp4_r_v_b_37')
// (9, 18, 'local_g0_0')
// (9, 18, 'lutff_3/in_1')
// (9, 18, 'sp4_r_v_b_24')
// (9, 19, 'sp4_r_v_b_13')
// (9, 20, 'sp4_r_v_b_0')
// (10, 11, 'neigh_op_tnr_7')
// (10, 12, 'neigh_op_rgt_7')
// (10, 12, 'sp4_h_r_3')
// (10, 12, 'sp4_r_v_b_46')
// (10, 12, 'sp4_v_t_44')
// (10, 13, 'neigh_op_bnr_7')
// (10, 13, 'sp4_r_v_b_35')
// (10, 13, 'sp4_v_b_44')
// (10, 14, 'sp4_r_v_b_22')
// (10, 14, 'sp4_v_b_33')
// (10, 15, 'sp4_r_v_b_11')
// (10, 15, 'sp4_v_b_20')
// (10, 16, 'sp4_h_r_9')
// (10, 16, 'sp4_v_b_9')
// (10, 16, 'sp4_v_t_37')
// (10, 17, 'sp4_v_b_37')
// (10, 18, 'sp4_v_b_24')
// (10, 19, 'local_g1_5')
// (10, 19, 'lutff_7/in_3')
// (10, 19, 'sp4_r_v_b_46')
// (10, 19, 'sp4_v_b_13')
// (10, 20, 'local_g0_0')
// (10, 20, 'lutff_5/in_1')
// (10, 20, 'sp4_h_r_6')
// (10, 20, 'sp4_r_v_b_35')
// (10, 20, 'sp4_v_b_0')
// (10, 21, 'sp4_r_v_b_22')
// (10, 22, 'sp4_r_v_b_11')
// (10, 23, 'local_g3_2')
// (10, 23, 'lutff_6/in_3')
// (10, 23, 'sp4_r_v_b_42')
// (10, 24, 'sp4_r_v_b_31')
// (10, 25, 'sp4_r_v_b_18')
// (10, 26, 'sp4_r_v_b_7')
// (11, 7, 'sp12_h_r_1')
// (11, 7, 'sp12_v_t_22')
// (11, 8, 'sp12_v_b_22')
// (11, 9, 'sp12_v_b_21')
// (11, 10, 'sp12_v_b_18')
// (11, 11, 'neigh_op_top_7')
// (11, 11, 'sp12_v_b_17')
// (11, 11, 'sp4_v_t_46')
// (11, 12, 'lutff_7/out')
// (11, 12, 'sp12_v_b_14')
// (11, 12, 'sp4_h_r_14')
// (11, 12, 'sp4_r_v_b_47')
// (11, 12, 'sp4_v_b_46')
// (11, 13, 'local_g1_7')
// (11, 13, 'lutff_5/in_3')
// (11, 13, 'neigh_op_bot_7')
// (11, 13, 'sp12_v_b_13')
// (11, 13, 'sp4_r_v_b_34')
// (11, 13, 'sp4_v_b_35')
// (11, 14, 'sp12_v_b_10')
// (11, 14, 'sp4_r_v_b_23')
// (11, 14, 'sp4_v_b_22')
// (11, 15, 'sp12_v_b_9')
// (11, 15, 'sp4_h_r_11')
// (11, 15, 'sp4_r_v_b_10')
// (11, 15, 'sp4_v_b_11')
// (11, 16, 'sp12_v_b_6')
// (11, 16, 'sp4_h_r_20')
// (11, 16, 'sp4_r_v_b_36')
// (11, 17, 'sp12_v_b_5')
// (11, 17, 'sp4_r_v_b_25')
// (11, 18, 'sp12_v_b_2')
// (11, 18, 'sp4_h_r_4')
// (11, 18, 'sp4_r_v_b_12')
// (11, 18, 'sp4_v_t_46')
// (11, 19, 'sp12_v_b_1')
// (11, 19, 'sp12_v_t_22')
// (11, 19, 'sp4_r_v_b_1')
// (11, 19, 'sp4_v_b_46')
// (11, 20, 'sp12_v_b_22')
// (11, 20, 'sp4_h_r_19')
// (11, 20, 'sp4_v_b_35')
// (11, 21, 'sp12_v_b_21')
// (11, 21, 'sp4_v_b_22')
// (11, 22, 'sp12_v_b_18')
// (11, 22, 'sp4_h_r_11')
// (11, 22, 'sp4_v_b_11')
// (11, 22, 'sp4_v_t_42')
// (11, 23, 'sp12_v_b_17')
// (11, 23, 'sp4_v_b_42')
// (11, 24, 'sp12_v_b_14')
// (11, 24, 'sp4_v_b_31')
// (11, 25, 'sp12_v_b_13')
// (11, 25, 'sp4_v_b_18')
// (11, 26, 'sp12_v_b_10')
// (11, 26, 'sp4_v_b_7')
// (11, 27, 'sp12_v_b_9')
// (11, 28, 'sp12_v_b_6')
// (11, 29, 'sp12_v_b_5')
// (11, 30, 'sp12_v_b_2')
// (11, 31, 'sp12_h_r_1')
// (11, 31, 'sp12_v_b_1')
// (12, 7, 'sp12_h_r_2')
// (12, 11, 'neigh_op_tnl_7')
// (12, 11, 'sp4_h_r_10')
// (12, 11, 'sp4_v_t_47')
// (12, 12, 'neigh_op_lft_7')
// (12, 12, 'sp4_h_r_27')
// (12, 12, 'sp4_v_b_47')
// (12, 13, 'local_g3_7')
// (12, 13, 'lutff_7/in_3')
// (12, 13, 'neigh_op_bnl_7')
// (12, 13, 'sp4_v_b_34')
// (12, 14, 'sp4_v_b_23')
// (12, 15, 'sp4_h_r_10')
// (12, 15, 'sp4_h_r_22')
// (12, 15, 'sp4_v_b_10')
// (12, 15, 'sp4_v_t_36')
// (12, 16, 'sp4_h_r_33')
// (12, 16, 'sp4_v_b_36')
// (12, 17, 'sp4_v_b_25')
// (12, 18, 'sp4_h_r_17')
// (12, 18, 'sp4_v_b_12')
// (12, 19, 'local_g1_1')
// (12, 19, 'lutff_7/in_3')
// (12, 19, 'sp4_v_b_1')
// (12, 20, 'local_g2_6')
// (12, 20, 'lutff_7/in_3')
// (12, 20, 'sp4_h_r_30')
// (12, 22, 'sp4_h_r_22')
// (12, 31, 'sp12_h_r_2')
// (13, 7, 'sp12_h_r_5')
// (13, 11, 'sp4_h_r_23')
// (13, 12, 'sp4_h_r_38')
// (13, 15, 'sp4_h_r_23')
// (13, 15, 'sp4_h_r_35')
// (13, 16, 'local_g2_4')
// (13, 16, 'lutff_5/in_3')
// (13, 16, 'sp4_h_r_44')
// (13, 18, 'sp4_h_r_28')
// (13, 20, 'sp4_h_r_43')
// (13, 22, 'sp4_h_r_35')
// (13, 31, 'sp12_h_r_5')
// (14, 7, 'sp12_h_r_6')
// (14, 11, 'sp4_h_r_34')
// (14, 12, 'sp4_h_l_38')
// (14, 12, 'sp4_h_r_6')
// (14, 12, 'sp4_r_v_b_40')
// (14, 13, 'local_g1_5')
// (14, 13, 'lutff_7/in_3')
// (14, 13, 'sp4_r_v_b_29')
// (14, 14, 'local_g3_0')
// (14, 14, 'lutff_0/in_1')
// (14, 14, 'sp4_r_v_b_16')
// (14, 15, 'local_g3_6')
// (14, 15, 'lutff_4/in_3')
// (14, 15, 'sp4_h_r_34')
// (14, 15, 'sp4_h_r_46')
// (14, 15, 'sp4_r_v_b_41')
// (14, 15, 'sp4_r_v_b_5')
// (14, 16, 'sp4_h_l_44')
// (14, 16, 'sp4_r_v_b_28')
// (14, 16, 'sp4_r_v_b_46')
// (14, 17, 'sp4_r_v_b_17')
// (14, 17, 'sp4_r_v_b_35')
// (14, 18, 'sp4_h_r_41')
// (14, 18, 'sp4_r_v_b_22')
// (14, 18, 'sp4_r_v_b_4')
// (14, 19, 'sp4_r_v_b_11')
// (14, 20, 'sp4_h_l_43')
// (14, 22, 'local_g2_6')
// (14, 22, 'lutff_5/in_3')
// (14, 22, 'sp4_h_r_46')
// (14, 31, 'sp12_h_r_6')
// (15, 7, 'sp12_h_r_9')
// (15, 7, 'sp4_h_r_4')
// (15, 8, 'sp4_r_v_b_41')
// (15, 9, 'sp4_r_v_b_28')
// (15, 10, 'sp4_r_v_b_17')
// (15, 11, 'sp4_h_r_10')
// (15, 11, 'sp4_h_r_47')
// (15, 11, 'sp4_r_v_b_4')
// (15, 11, 'sp4_v_t_40')
// (15, 12, 'sp4_h_r_19')
// (15, 12, 'sp4_v_b_40')
// (15, 13, 'sp4_v_b_29')
// (15, 14, 'sp4_v_b_16')
// (15, 14, 'sp4_v_t_41')
// (15, 15, 'local_g3_7')
// (15, 15, 'lutff_7/in_3')
// (15, 15, 'sp4_h_l_46')
// (15, 15, 'sp4_h_r_47')
// (15, 15, 'sp4_v_b_41')
// (15, 15, 'sp4_v_b_5')
// (15, 15, 'sp4_v_t_46')
// (15, 16, 'sp4_r_v_b_38')
// (15, 16, 'sp4_v_b_28')
// (15, 16, 'sp4_v_b_46')
// (15, 17, 'local_g1_1')
// (15, 17, 'lutff_7/in_3')
// (15, 17, 'sp4_r_v_b_27')
// (15, 17, 'sp4_v_b_17')
// (15, 17, 'sp4_v_b_35')
// (15, 18, 'local_g0_4')
// (15, 18, 'lutff_7/in_3')
// (15, 18, 'sp4_h_l_41')
// (15, 18, 'sp4_r_v_b_14')
// (15, 18, 'sp4_v_b_22')
// (15, 18, 'sp4_v_b_4')
// (15, 19, 'local_g1_3')
// (15, 19, 'lutff_7/in_3')
// (15, 19, 'sp4_r_v_b_3')
// (15, 19, 'sp4_v_b_11')
// (15, 20, 'sp4_r_v_b_38')
// (15, 21, 'sp4_r_v_b_27')
// (15, 22, 'sp4_h_l_46')
// (15, 22, 'sp4_r_v_b_14')
// (15, 23, 'sp4_r_v_b_3')
// (15, 31, 'sp12_h_r_9')
// (16, 7, 'sp12_h_r_10')
// (16, 7, 'sp4_h_r_17')
// (16, 7, 'sp4_v_t_41')
// (16, 8, 'sp4_v_b_41')
// (16, 9, 'local_g2_4')
// (16, 9, 'lutff_1/in_3')
// (16, 9, 'sp4_v_b_28')
// (16, 10, 'sp4_v_b_17')
// (16, 11, 'local_g1_7')
// (16, 11, 'lutff_7/in_3')
// (16, 11, 'sp4_h_l_47')
// (16, 11, 'sp4_h_r_23')
// (16, 11, 'sp4_v_b_4')
// (16, 12, 'sp4_h_r_30')
// (16, 15, 'sp4_h_l_47')
// (16, 15, 'sp4_v_t_38')
// (16, 16, 'local_g3_6')
// (16, 16, 'lutff_7/in_0')
// (16, 16, 'sp4_v_b_38')
// (16, 17, 'local_g3_3')
// (16, 17, 'lutff_7/in_3')
// (16, 17, 'sp4_v_b_27')
// (16, 18, 'local_g0_6')
// (16, 18, 'lutff_7/in_3')
// (16, 18, 'sp4_v_b_14')
// (16, 19, 'local_g1_3')
// (16, 19, 'lutff_5/in_3')
// (16, 19, 'sp4_h_r_9')
// (16, 19, 'sp4_v_b_3')
// (16, 19, 'sp4_v_t_38')
// (16, 20, 'sp4_v_b_38')
// (16, 21, 'local_g2_3')
// (16, 21, 'lutff_5/in_0')
// (16, 21, 'sp4_v_b_27')
// (16, 22, 'sp4_v_b_14')
// (16, 23, 'sp4_v_b_3')
// (16, 31, 'sp12_h_r_10')
// (17, 7, 'sp12_h_r_13')
// (17, 7, 'sp4_h_r_28')
// (17, 7, 'sp4_h_r_6')
// (17, 11, 'sp4_h_r_34')
// (17, 12, 'sp4_h_r_43')
// (17, 13, 'sp4_r_v_b_46')
// (17, 14, 'sp4_r_v_b_35')
// (17, 15, 'sp4_r_v_b_22')
// (17, 16, 'sp4_r_v_b_11')
// (17, 17, 'sp4_r_v_b_46')
// (17, 18, 'sp4_r_v_b_35')
// (17, 19, 'sp4_h_r_20')
// (17, 19, 'sp4_r_v_b_22')
// (17, 20, 'sp4_r_v_b_11')
// (17, 21, 'sp4_r_v_b_39')
// (17, 22, 'sp4_r_v_b_26')
// (17, 23, 'sp4_r_v_b_15')
// (17, 24, 'sp4_r_v_b_2')
// (17, 31, 'sp12_h_r_13')
// (17, 31, 'sp4_h_r_6')
// (18, 7, 'sp12_h_r_14')
// (18, 7, 'sp4_h_r_19')
// (18, 7, 'sp4_h_r_41')
// (18, 8, 'sp4_r_v_b_44')
// (18, 9, 'sp4_r_v_b_33')
// (18, 10, 'sp4_r_v_b_20')
// (18, 11, 'local_g3_7')
// (18, 11, 'lutff_3/in_3')
// (18, 11, 'sp4_h_r_47')
// (18, 11, 'sp4_r_v_b_9')
// (18, 12, 'local_g0_1')
// (18, 12, 'lutff_7/in_0')
// (18, 12, 'sp4_h_l_43')
// (18, 12, 'sp4_h_r_9')
// (18, 12, 'sp4_v_t_46')
// (18, 13, 'sp4_v_b_46')
// (18, 14, 'sp4_v_b_35')
// (18, 15, 'sp4_v_b_22')
// (18, 16, 'sp4_h_r_5')
// (18, 16, 'sp4_v_b_11')
// (18, 16, 'sp4_v_t_46')
// (18, 17, 'local_g2_6')
// (18, 17, 'lutff_3/in_3')
// (18, 17, 'sp4_v_b_46')
// (18, 18, 'sp4_v_b_35')
// (18, 19, 'sp4_h_r_33')
// (18, 19, 'sp4_v_b_22')
// (18, 20, 'sp4_h_r_5')
// (18, 20, 'sp4_v_b_11')
// (18, 20, 'sp4_v_t_39')
// (18, 21, 'sp4_v_b_39')
// (18, 22, 'sp4_v_b_26')
// (18, 23, 'sp4_v_b_15')
// (18, 24, 'local_g1_2')
// (18, 24, 'lutff_6/in_3')
// (18, 24, 'sp4_v_b_2')
// (18, 31, 'sp12_h_r_14')
// (18, 31, 'sp4_h_r_19')
// (19, 7, 'sp12_h_r_17')
// (19, 7, 'sp4_h_l_41')
// (19, 7, 'sp4_h_r_30')
// (19, 7, 'sp4_v_t_44')
// (19, 8, 'sp4_v_b_44')
// (19, 9, 'local_g2_1')
// (19, 9, 'lutff_0/in_3')
// (19, 9, 'sp4_v_b_33')
// (19, 10, 'local_g0_4')
// (19, 10, 'lutff_7/in_3')
// (19, 10, 'sp4_v_b_20')
// (19, 11, 'local_g0_1')
// (19, 11, 'lutff_7/in_0')
// (19, 11, 'sp4_h_l_47')
// (19, 11, 'sp4_v_b_9')
// (19, 12, 'sp4_h_r_20')
// (19, 16, 'local_g0_0')
// (19, 16, 'lutff_7/in_1')
// (19, 16, 'sp4_h_r_16')
// (19, 19, 'local_g3_4')
// (19, 19, 'lutff_6/in_3')
// (19, 19, 'sp4_h_r_44')
// (19, 20, 'sp4_h_r_16')
// (19, 31, 'sp12_h_r_17')
// (19, 31, 'sp4_h_r_30')
// (20, 7, 'sp12_h_r_18')
// (20, 7, 'sp4_h_r_43')
// (20, 8, 'sp4_r_v_b_43')
// (20, 9, 'sp4_r_v_b_30')
// (20, 10, 'sp4_r_v_b_19')
// (20, 11, 'local_g1_6')
// (20, 11, 'lutff_6/in_3')
// (20, 11, 'sp4_r_v_b_6')
// (20, 12, 'local_g3_1')
// (20, 12, 'lutff_7/in_3')
// (20, 12, 'sp4_h_r_33')
// (20, 16, 'local_g3_5')
// (20, 16, 'lutff_7/in_3')
// (20, 16, 'sp4_h_r_29')
// (20, 19, 'local_g1_5')
// (20, 19, 'lutff_7/in_3')
// (20, 19, 'sp4_h_l_44')
// (20, 19, 'sp4_h_r_5')
// (20, 20, 'local_g3_5')
// (20, 20, 'lutff_7/in_3')
// (20, 20, 'sp4_h_r_29')
// (20, 24, 'sp4_r_v_b_43')
// (20, 25, 'local_g0_6')
// (20, 25, 'lutff_7/in_3')
// (20, 25, 'sp4_r_v_b_30')
// (20, 26, 'sp4_r_v_b_19')
// (20, 27, 'sp4_r_v_b_6')
// (20, 28, 'sp4_r_v_b_43')
// (20, 29, 'sp4_r_v_b_30')
// (20, 30, 'sp4_r_v_b_19')
// (20, 31, 'sp12_h_r_18')
// (20, 31, 'sp4_h_r_43')
// (20, 31, 'sp4_r_v_b_6')
// (21, 7, 'sp12_h_r_21')
// (21, 7, 'sp4_h_l_43')
// (21, 7, 'sp4_h_r_10')
// (21, 7, 'sp4_v_t_43')
// (21, 8, 'sp4_v_b_43')
// (21, 9, 'sp4_v_b_30')
// (21, 10, 'sp4_v_b_19')
// (21, 11, 'local_g0_6')
// (21, 11, 'lutff_7/in_3')
// (21, 11, 'sp4_v_b_6')
// (21, 12, 'local_g3_4')
// (21, 12, 'lutff_7/in_0')
// (21, 12, 'sp4_h_r_44')
// (21, 13, 'sp4_r_v_b_44')
// (21, 14, 'sp4_r_v_b_33')
// (21, 15, 'sp4_r_v_b_20')
// (21, 16, 'sp4_h_r_40')
// (21, 16, 'sp4_r_v_b_9')
// (21, 19, 'sp4_h_r_16')
// (21, 20, 'local_g2_0')
// (21, 20, 'lutff_7/in_3')
// (21, 20, 'sp4_h_r_40')
// (21, 21, 'sp4_r_v_b_47')
// (21, 22, 'sp4_r_v_b_34')
// (21, 23, 'sp4_r_v_b_23')
// (21, 23, 'sp4_v_t_43')
// (21, 24, 'sp4_r_v_b_10')
// (21, 24, 'sp4_v_b_43')
// (21, 25, 'sp4_v_b_30')
// (21, 26, 'sp4_v_b_19')
// (21, 27, 'sp4_v_b_6')
// (21, 27, 'sp4_v_t_43')
// (21, 28, 'sp4_v_b_43')
// (21, 29, 'sp4_v_b_30')
// (21, 30, 'sp4_v_b_19')
// (21, 31, 'sp12_h_r_21')
// (21, 31, 'sp4_h_l_43')
// (21, 31, 'sp4_v_b_6')
// (22, 7, 'sp12_h_r_22')
// (22, 7, 'sp4_h_r_23')
// (22, 12, 'local_g1_1')
// (22, 12, 'lutff_7/in_3')
// (22, 12, 'sp4_h_l_44')
// (22, 12, 'sp4_h_r_9')
// (22, 12, 'sp4_v_t_44')
// (22, 13, 'sp4_v_b_44')
// (22, 14, 'local_g3_1')
// (22, 14, 'lutff_7/in_3')
// (22, 14, 'sp4_v_b_33')
// (22, 15, 'sp4_v_b_20')
// (22, 16, 'sp4_h_l_40')
// (22, 16, 'sp4_h_r_1')
// (22, 16, 'sp4_v_b_9')
// (22, 19, 'sp4_h_r_29')
// (22, 20, 'sp4_h_l_40')
// (22, 20, 'sp4_h_r_1')
// (22, 20, 'sp4_v_t_47')
// (22, 21, 'local_g3_7')
// (22, 21, 'lutff_7/in_3')
// (22, 21, 'sp4_v_b_47')
// (22, 22, 'sp4_v_b_34')
// (22, 23, 'local_g1_7')
// (22, 23, 'lutff_7/in_3')
// (22, 23, 'sp4_v_b_23')
// (22, 24, 'local_g0_2')
// (22, 24, 'lutff_1/in_3')
// (22, 24, 'sp4_v_b_10')
// (22, 31, 'sp12_h_r_22')
// (23, 7, 'sp12_h_l_22')
// (23, 7, 'sp12_v_t_22')
// (23, 7, 'sp4_h_r_34')
// (23, 8, 'sp12_v_b_22')
// (23, 9, 'sp12_v_b_21')
// (23, 10, 'sp12_v_b_18')
// (23, 11, 'sp12_v_b_17')
// (23, 12, 'local_g0_4')
// (23, 12, 'lutff_7/in_3')
// (23, 12, 'sp12_v_b_14')
// (23, 12, 'sp4_h_r_20')
// (23, 13, 'sp12_v_b_13')
// (23, 14, 'local_g3_2')
// (23, 14, 'lutff_7/in_0')
// (23, 14, 'sp12_v_b_10')
// (23, 15, 'local_g3_1')
// (23, 15, 'lutff_7/in_3')
// (23, 15, 'sp12_v_b_9')
// (23, 16, 'local_g0_4')
// (23, 16, 'lutff_7/in_3')
// (23, 16, 'sp12_v_b_6')
// (23, 16, 'sp4_h_r_12')
// (23, 17, 'sp12_v_b_5')
// (23, 18, 'sp12_v_b_2')
// (23, 19, 'sp12_v_b_1')
// (23, 19, 'sp12_v_t_22')
// (23, 19, 'sp4_h_r_40')
// (23, 20, 'local_g0_4')
// (23, 20, 'lutff_7/in_3')
// (23, 20, 'sp12_v_b_22')
// (23, 20, 'sp4_h_r_12')
// (23, 21, 'sp12_v_b_21')
// (23, 22, 'local_g2_2')
// (23, 22, 'lutff_5/in_3')
// (23, 22, 'sp12_v_b_18')
// (23, 23, 'sp12_v_b_17')
// (23, 24, 'sp12_v_b_14')
// (23, 25, 'sp12_v_b_13')
// (23, 26, 'sp12_v_b_10')
// (23, 27, 'sp12_v_b_9')
// (23, 28, 'sp12_v_b_6')
// (23, 29, 'sp12_v_b_5')
// (23, 30, 'sp12_v_b_2')
// (23, 31, 'sp12_h_l_22')
// (23, 31, 'sp12_v_b_1')
// (24, 7, 'sp4_h_r_47')
// (24, 8, 'sp4_r_v_b_38')
// (24, 9, 'sp4_r_v_b_27')
// (24, 10, 'sp4_r_v_b_14')
// (24, 11, 'sp4_r_v_b_3')
// (24, 12, 'sp4_h_r_33')
// (24, 12, 'sp4_r_v_b_43')
// (24, 12, 'sp4_r_v_b_46')
// (24, 13, 'local_g2_3')
// (24, 13, 'lutff_2/in_3')
// (24, 13, 'sp4_r_v_b_30')
// (24, 13, 'sp4_r_v_b_35')
// (24, 14, 'local_g3_3')
// (24, 14, 'lutff_7/in_3')
// (24, 14, 'sp4_r_v_b_19')
// (24, 14, 'sp4_r_v_b_22')
// (24, 15, 'local_g1_6')
// (24, 15, 'lutff_3/in_0')
// (24, 15, 'sp4_r_v_b_11')
// (24, 15, 'sp4_r_v_b_6')
// (24, 16, 'local_g2_1')
// (24, 16, 'lutff_2/in_3')
// (24, 16, 'sp4_h_r_25')
// (24, 16, 'sp4_r_v_b_43')
// (24, 17, 'local_g0_6')
// (24, 17, 'lutff_7/in_3')
// (24, 17, 'sp4_r_v_b_30')
// (24, 18, 'sp4_r_v_b_19')
// (24, 19, 'sp4_h_l_40')
// (24, 19, 'sp4_r_v_b_6')
// (24, 20, 'sp4_h_r_25')
// (25, 7, 'sp4_h_l_47')
// (25, 7, 'sp4_v_t_38')
// (25, 8, 'sp4_v_b_38')
// (25, 9, 'sp4_v_b_27')
// (25, 10, 'sp4_v_b_14')
// (25, 11, 'sp4_v_b_3')
// (25, 11, 'sp4_v_t_43')
// (25, 11, 'sp4_v_t_46')
// (25, 12, 'sp4_h_r_44')
// (25, 12, 'sp4_v_b_43')
// (25, 12, 'sp4_v_b_46')
// (25, 13, 'sp4_v_b_30')
// (25, 13, 'sp4_v_b_35')
// (25, 14, 'sp4_v_b_19')
// (25, 14, 'sp4_v_b_22')
// (25, 15, 'sp4_v_b_11')
// (25, 15, 'sp4_v_b_6')
// (25, 15, 'sp4_v_t_43')
// (25, 16, 'sp4_h_r_36')
// (25, 16, 'sp4_v_b_43')
// (25, 17, 'sp4_v_b_30')
// (25, 18, 'sp4_v_b_19')
// (25, 19, 'sp4_v_b_6')
// (25, 20, 'sp4_h_r_36')
// (26, 12, 'sp4_h_l_44')
// (26, 16, 'sp4_h_l_36')
// (26, 20, 'sp4_h_l_36')

wire n219;
// (9, 14, 'neigh_op_tnr_0')
// (9, 15, 'local_g2_0')
// (9, 15, 'lutff_1/in_3')
// (9, 15, 'neigh_op_rgt_0')
// (9, 16, 'neigh_op_bnr_0')
// (10, 14, 'neigh_op_top_0')
// (10, 15, 'lutff_0/out')
// (10, 16, 'neigh_op_bot_0')
// (11, 14, 'neigh_op_tnl_0')
// (11, 15, 'neigh_op_lft_0')
// (11, 16, 'neigh_op_bnl_0')

reg n220 = 0;
// (9, 14, 'neigh_op_tnr_1')
// (9, 15, 'local_g2_1')
// (9, 15, 'lutff_4/in_3')
// (9, 15, 'neigh_op_rgt_1')
// (9, 16, 'neigh_op_bnr_1')
// (10, 14, 'neigh_op_top_1')
// (10, 15, 'local_g3_1')
// (10, 15, 'lutff_1/in_1')
// (10, 15, 'lutff_1/out')
// (10, 16, 'neigh_op_bot_1')
// (11, 14, 'neigh_op_tnl_1')
// (11, 15, 'neigh_op_lft_1')
// (11, 16, 'neigh_op_bnl_1')

reg n221 = 0;
// (9, 14, 'neigh_op_tnr_2')
// (9, 15, 'local_g3_2')
// (9, 15, 'lutff_4/in_1')
// (9, 15, 'neigh_op_rgt_2')
// (9, 16, 'neigh_op_bnr_2')
// (10, 14, 'neigh_op_top_2')
// (10, 15, 'local_g1_2')
// (10, 15, 'lutff_2/in_1')
// (10, 15, 'lutff_2/out')
// (10, 16, 'neigh_op_bot_2')
// (11, 14, 'neigh_op_tnl_2')
// (11, 15, 'neigh_op_lft_2')
// (11, 16, 'neigh_op_bnl_2')

reg n222 = 0;
// (9, 14, 'neigh_op_tnr_3')
// (9, 15, 'local_g3_3')
// (9, 15, 'lutff_4/in_0')
// (9, 15, 'neigh_op_rgt_3')
// (9, 16, 'neigh_op_bnr_3')
// (10, 14, 'neigh_op_top_3')
// (10, 15, 'local_g1_3')
// (10, 15, 'lutff_3/in_1')
// (10, 15, 'lutff_3/out')
// (10, 16, 'neigh_op_bot_3')
// (11, 14, 'neigh_op_tnl_3')
// (11, 15, 'neigh_op_lft_3')
// (11, 16, 'neigh_op_bnl_3')

reg n223 = 0;
// (9, 14, 'neigh_op_tnr_4')
// (9, 15, 'local_g2_4')
// (9, 15, 'lutff_4/in_2')
// (9, 15, 'neigh_op_rgt_4')
// (9, 16, 'neigh_op_bnr_4')
// (10, 14, 'neigh_op_top_4')
// (10, 15, 'local_g3_4')
// (10, 15, 'lutff_4/in_1')
// (10, 15, 'lutff_4/out')
// (10, 16, 'neigh_op_bot_4')
// (11, 14, 'neigh_op_tnl_4')
// (11, 15, 'neigh_op_lft_4')
// (11, 16, 'neigh_op_bnl_4')

reg n224 = 0;
// (9, 14, 'neigh_op_tnr_5')
// (9, 15, 'local_g2_5')
// (9, 15, 'lutff_7/in_0')
// (9, 15, 'neigh_op_rgt_5')
// (9, 16, 'neigh_op_bnr_5')
// (10, 14, 'neigh_op_top_5')
// (10, 15, 'local_g1_5')
// (10, 15, 'lutff_5/in_1')
// (10, 15, 'lutff_5/out')
// (10, 16, 'neigh_op_bot_5')
// (11, 14, 'neigh_op_tnl_5')
// (11, 15, 'neigh_op_lft_5')
// (11, 16, 'neigh_op_bnl_5')

reg n225 = 0;
// (9, 14, 'neigh_op_tnr_6')
// (9, 15, 'local_g2_6')
// (9, 15, 'lutff_7/in_3')
// (9, 15, 'neigh_op_rgt_6')
// (9, 16, 'neigh_op_bnr_6')
// (10, 14, 'neigh_op_top_6')
// (10, 15, 'local_g1_6')
// (10, 15, 'lutff_6/in_1')
// (10, 15, 'lutff_6/out')
// (10, 16, 'neigh_op_bot_6')
// (11, 14, 'neigh_op_tnl_6')
// (11, 15, 'neigh_op_lft_6')
// (11, 16, 'neigh_op_bnl_6')

reg n226 = 0;
// (9, 14, 'neigh_op_tnr_7')
// (9, 15, 'local_g3_7')
// (9, 15, 'lutff_7/in_1')
// (9, 15, 'neigh_op_rgt_7')
// (9, 16, 'neigh_op_bnr_7')
// (10, 14, 'neigh_op_top_7')
// (10, 15, 'local_g3_7')
// (10, 15, 'lutff_7/in_1')
// (10, 15, 'lutff_7/out')
// (10, 16, 'neigh_op_bot_7')
// (11, 14, 'neigh_op_tnl_7')
// (11, 15, 'neigh_op_lft_7')
// (11, 16, 'neigh_op_bnl_7')

reg n227 = 0;
// (9, 14, 'sp4_r_v_b_45')
// (9, 15, 'local_g0_3')
// (9, 15, 'lutff_1/in_0')
// (9, 15, 'sp4_r_v_b_32')
// (9, 16, 'neigh_op_tnr_4')
// (9, 16, 'sp4_r_v_b_21')
// (9, 17, 'neigh_op_rgt_4')
// (9, 17, 'sp4_r_v_b_8')
// (9, 18, 'neigh_op_bnr_4')
// (10, 13, 'sp4_v_t_45')
// (10, 14, 'sp4_v_b_45')
// (10, 15, 'sp4_v_b_32')
// (10, 16, 'neigh_op_top_4')
// (10, 16, 'sp4_v_b_21')
// (10, 17, 'local_g3_4')
// (10, 17, 'lutff_4/in_1')
// (10, 17, 'lutff_4/out')
// (10, 17, 'sp4_v_b_8')
// (10, 18, 'neigh_op_bot_4')
// (11, 16, 'neigh_op_tnl_4')
// (11, 17, 'neigh_op_lft_4')
// (11, 18, 'neigh_op_bnl_4')

reg n228 = 0;
// (9, 14, 'sp4_r_v_b_47')
// (9, 15, 'local_g0_1')
// (9, 15, 'lutff_1/in_2')
// (9, 15, 'sp4_r_v_b_34')
// (9, 16, 'neigh_op_tnr_5')
// (9, 16, 'sp4_r_v_b_23')
// (9, 17, 'neigh_op_rgt_5')
// (9, 17, 'sp4_r_v_b_10')
// (9, 18, 'neigh_op_bnr_5')
// (10, 13, 'sp4_v_t_47')
// (10, 14, 'sp4_v_b_47')
// (10, 15, 'sp4_v_b_34')
// (10, 16, 'neigh_op_top_5')
// (10, 16, 'sp4_v_b_23')
// (10, 17, 'local_g1_5')
// (10, 17, 'lutff_5/in_1')
// (10, 17, 'lutff_5/out')
// (10, 17, 'sp4_v_b_10')
// (10, 18, 'neigh_op_bot_5')
// (11, 16, 'neigh_op_tnl_5')
// (11, 17, 'neigh_op_lft_5')
// (11, 18, 'neigh_op_bnl_5')

reg n229 = 0;
// (9, 15, 'local_g3_0')
// (9, 15, 'lutff_7/in_2')
// (9, 15, 'neigh_op_tnr_0')
// (9, 16, 'neigh_op_rgt_0')
// (9, 17, 'neigh_op_bnr_0')
// (10, 15, 'neigh_op_top_0')
// (10, 16, 'local_g3_0')
// (10, 16, 'lutff_0/in_1')
// (10, 16, 'lutff_0/out')
// (10, 17, 'neigh_op_bot_0')
// (11, 15, 'neigh_op_tnl_0')
// (11, 16, 'neigh_op_lft_0')
// (11, 17, 'neigh_op_bnl_0')

wire n230;
// (9, 15, 'lutff_5/lout')
// (9, 15, 'lutff_6/in_2')

reg n231 = 0;
// (9, 15, 'neigh_op_tnr_1')
// (9, 16, 'local_g3_1')
// (9, 16, 'lutff_0/in_0')
// (9, 16, 'neigh_op_rgt_1')
// (9, 17, 'neigh_op_bnr_1')
// (10, 15, 'neigh_op_top_1')
// (10, 16, 'local_g3_1')
// (10, 16, 'lutff_1/in_1')
// (10, 16, 'lutff_1/out')
// (10, 17, 'neigh_op_bot_1')
// (11, 15, 'neigh_op_tnl_1')
// (11, 16, 'neigh_op_lft_1')
// (11, 17, 'neigh_op_bnl_1')

reg n232 = 0;
// (9, 15, 'neigh_op_tnr_2')
// (9, 16, 'local_g3_2')
// (9, 16, 'lutff_0/in_3')
// (9, 16, 'neigh_op_rgt_2')
// (9, 17, 'neigh_op_bnr_2')
// (10, 15, 'neigh_op_top_2')
// (10, 16, 'local_g1_2')
// (10, 16, 'lutff_2/in_1')
// (10, 16, 'lutff_2/out')
// (10, 17, 'neigh_op_bot_2')
// (11, 15, 'neigh_op_tnl_2')
// (11, 16, 'neigh_op_lft_2')
// (11, 17, 'neigh_op_bnl_2')

reg n233 = 0;
// (9, 15, 'neigh_op_tnr_3')
// (9, 16, 'local_g2_3')
// (9, 16, 'lutff_0/in_1')
// (9, 16, 'neigh_op_rgt_3')
// (9, 17, 'neigh_op_bnr_3')
// (10, 15, 'neigh_op_top_3')
// (10, 16, 'local_g1_3')
// (10, 16, 'lutff_3/in_1')
// (10, 16, 'lutff_3/out')
// (10, 17, 'neigh_op_bot_3')
// (11, 15, 'neigh_op_tnl_3')
// (11, 16, 'neigh_op_lft_3')
// (11, 17, 'neigh_op_bnl_3')

reg n234 = 0;
// (9, 15, 'neigh_op_tnr_4')
// (9, 16, 'local_g2_4')
// (9, 16, 'lutff_0/in_2')
// (9, 16, 'neigh_op_rgt_4')
// (9, 17, 'neigh_op_bnr_4')
// (10, 15, 'neigh_op_top_4')
// (10, 16, 'local_g3_4')
// (10, 16, 'lutff_4/in_1')
// (10, 16, 'lutff_4/out')
// (10, 17, 'neigh_op_bot_4')
// (11, 15, 'neigh_op_tnl_4')
// (11, 16, 'neigh_op_lft_4')
// (11, 17, 'neigh_op_bnl_4')

reg n235 = 0;
// (9, 15, 'neigh_op_tnr_5')
// (9, 16, 'local_g2_5')
// (9, 16, 'lutff_2/in_3')
// (9, 16, 'neigh_op_rgt_5')
// (9, 17, 'neigh_op_bnr_5')
// (10, 15, 'neigh_op_top_5')
// (10, 16, 'local_g1_5')
// (10, 16, 'lutff_5/in_1')
// (10, 16, 'lutff_5/out')
// (10, 17, 'neigh_op_bot_5')
// (11, 15, 'neigh_op_tnl_5')
// (11, 16, 'neigh_op_lft_5')
// (11, 17, 'neigh_op_bnl_5')

reg n236 = 0;
// (9, 15, 'neigh_op_tnr_6')
// (9, 16, 'local_g3_6')
// (9, 16, 'lutff_2/in_1')
// (9, 16, 'neigh_op_rgt_6')
// (9, 17, 'neigh_op_bnr_6')
// (10, 15, 'neigh_op_top_6')
// (10, 16, 'local_g1_6')
// (10, 16, 'lutff_6/in_1')
// (10, 16, 'lutff_6/out')
// (10, 17, 'neigh_op_bot_6')
// (11, 15, 'neigh_op_tnl_6')
// (11, 16, 'neigh_op_lft_6')
// (11, 17, 'neigh_op_bnl_6')

reg n237 = 0;
// (9, 15, 'neigh_op_tnr_7')
// (9, 16, 'local_g3_7')
// (9, 16, 'lutff_2/in_0')
// (9, 16, 'neigh_op_rgt_7')
// (9, 17, 'neigh_op_bnr_7')
// (10, 15, 'neigh_op_top_7')
// (10, 16, 'local_g3_7')
// (10, 16, 'lutff_7/in_1')
// (10, 16, 'lutff_7/out')
// (10, 17, 'neigh_op_bot_7')
// (11, 15, 'neigh_op_tnl_7')
// (11, 16, 'neigh_op_lft_7')
// (11, 17, 'neigh_op_bnl_7')

wire n238;
// (9, 15, 'sp12_h_r_1')
// (10, 15, 'sp12_h_r_2')
// (11, 15, 'sp12_h_r_5')
// (12, 15, 'sp12_h_r_6')
// (13, 15, 'sp12_h_r_9')
// (14, 15, 'sp12_h_r_10')
// (15, 14, 'neigh_op_tnr_3')
// (15, 15, 'neigh_op_rgt_3')
// (15, 15, 'sp12_h_r_13')
// (15, 15, 'sp4_h_r_11')
// (15, 16, 'local_g1_3')
// (15, 16, 'lutff_1/in_3')
// (15, 16, 'neigh_op_bnr_3')
// (16, 14, 'neigh_op_top_3')
// (16, 14, 'sp12_v_t_22')
// (16, 15, 'lutff_3/out')
// (16, 15, 'sp12_h_r_14')
// (16, 15, 'sp12_v_b_22')
// (16, 15, 'sp4_h_r_22')
// (16, 16, 'neigh_op_bot_3')
// (16, 16, 'sp12_v_b_21')
// (16, 17, 'sp12_v_b_18')
// (16, 18, 'sp12_v_b_17')
// (16, 19, 'sp12_v_b_14')
// (16, 20, 'local_g3_5')
// (16, 20, 'lutff_1/in_3')
// (16, 20, 'lutff_2/in_0')
// (16, 20, 'lutff_3/in_3')
// (16, 20, 'lutff_7/in_3')
// (16, 20, 'sp12_v_b_13')
// (16, 21, 'sp12_v_b_10')
// (16, 22, 'sp12_v_b_9')
// (16, 23, 'sp12_v_b_6')
// (16, 24, 'sp12_v_b_5')
// (16, 25, 'sp12_v_b_2')
// (16, 26, 'sp12_v_b_1')
// (17, 14, 'neigh_op_tnl_3')
// (17, 15, 'neigh_op_lft_3')
// (17, 15, 'sp12_h_r_17')
// (17, 15, 'sp4_h_r_35')
// (17, 16, 'neigh_op_bnl_3')
// (18, 15, 'sp12_h_r_18')
// (18, 15, 'sp4_h_r_46')
// (19, 15, 'sp12_h_r_21')
// (19, 15, 'sp4_h_l_46')
// (19, 15, 'sp4_h_r_11')
// (20, 15, 'local_g0_6')
// (20, 15, 'lutff_0/in_0')
// (20, 15, 'lutff_1/in_3')
// (20, 15, 'lutff_3/in_3')
// (20, 15, 'lutff_5/in_3')
// (20, 15, 'sp12_h_r_22')
// (20, 15, 'sp4_h_r_22')
// (21, 15, 'sp12_h_l_22')
// (21, 15, 'sp4_h_r_35')
// (22, 15, 'local_g3_6')
// (22, 15, 'lutff_1/in_0')
// (22, 15, 'lutff_2/in_3')
// (22, 15, 'lutff_3/in_0')
// (22, 15, 'lutff_6/in_3')
// (22, 15, 'lutff_7/in_0')
// (22, 15, 'sp4_h_r_46')
// (23, 15, 'sp4_h_l_46')

reg n239 = 0;
// (9, 15, 'sp4_r_v_b_37')
// (9, 16, 'local_g0_0')
// (9, 16, 'lutff_2/in_2')
// (9, 16, 'sp4_r_v_b_24')
// (9, 17, 'neigh_op_tnr_0')
// (9, 17, 'sp4_r_v_b_13')
// (9, 18, 'neigh_op_rgt_0')
// (9, 18, 'sp4_r_v_b_0')
// (9, 19, 'neigh_op_bnr_0')
// (10, 14, 'sp4_v_t_37')
// (10, 15, 'sp4_v_b_37')
// (10, 16, 'sp4_v_b_24')
// (10, 17, 'neigh_op_top_0')
// (10, 17, 'sp4_v_b_13')
// (10, 18, 'local_g1_0')
// (10, 18, 'lutff_0/in_1')
// (10, 18, 'lutff_0/out')
// (10, 18, 'sp4_v_b_0')
// (10, 19, 'neigh_op_bot_0')
// (11, 17, 'neigh_op_tnl_0')
// (11, 18, 'neigh_op_lft_0')
// (11, 19, 'neigh_op_bnl_0')

reg n240 = 0;
// (9, 15, 'sp4_r_v_b_42')
// (9, 16, 'local_g0_7')
// (9, 16, 'lutff_1/in_0')
// (9, 16, 'neigh_op_tnr_1')
// (9, 16, 'sp4_r_v_b_31')
// (9, 17, 'neigh_op_rgt_1')
// (9, 17, 'sp4_r_v_b_18')
// (9, 18, 'neigh_op_bnr_1')
// (9, 18, 'sp4_r_v_b_7')
// (10, 14, 'sp4_v_t_42')
// (10, 15, 'sp4_v_b_42')
// (10, 16, 'neigh_op_top_1')
// (10, 16, 'sp4_v_b_31')
// (10, 17, 'local_g3_1')
// (10, 17, 'lutff_1/in_1')
// (10, 17, 'lutff_1/out')
// (10, 17, 'sp4_v_b_18')
// (10, 18, 'neigh_op_bot_1')
// (10, 18, 'sp4_v_b_7')
// (11, 16, 'neigh_op_tnl_1')
// (11, 17, 'neigh_op_lft_1')
// (11, 18, 'neigh_op_bnl_1')

reg n241 = 0;
// (9, 16, 'local_g2_2')
// (9, 16, 'lutff_1/in_3')
// (9, 16, 'neigh_op_tnr_2')
// (9, 17, 'neigh_op_rgt_2')
// (9, 18, 'neigh_op_bnr_2')
// (10, 16, 'neigh_op_top_2')
// (10, 17, 'local_g1_2')
// (10, 17, 'lutff_2/in_1')
// (10, 17, 'lutff_2/out')
// (10, 18, 'neigh_op_bot_2')
// (11, 16, 'neigh_op_tnl_2')
// (11, 17, 'neigh_op_lft_2')
// (11, 18, 'neigh_op_bnl_2')

reg n242 = 0;
// (9, 16, 'local_g3_0')
// (9, 16, 'lutff_1/in_2')
// (9, 16, 'neigh_op_tnr_0')
// (9, 17, 'neigh_op_rgt_0')
// (9, 18, 'neigh_op_bnr_0')
// (10, 16, 'neigh_op_top_0')
// (10, 17, 'local_g3_0')
// (10, 17, 'lutff_0/in_1')
// (10, 17, 'lutff_0/out')
// (10, 18, 'neigh_op_bot_0')
// (11, 16, 'neigh_op_tnl_0')
// (11, 17, 'neigh_op_lft_0')
// (11, 18, 'neigh_op_bnl_0')

reg n243 = 0;
// (9, 16, 'local_g3_3')
// (9, 16, 'lutff_1/in_1')
// (9, 16, 'neigh_op_tnr_3')
// (9, 17, 'neigh_op_rgt_3')
// (9, 18, 'neigh_op_bnr_3')
// (10, 16, 'neigh_op_top_3')
// (10, 17, 'local_g1_3')
// (10, 17, 'lutff_3/in_1')
// (10, 17, 'lutff_3/out')
// (10, 18, 'neigh_op_bot_3')
// (11, 16, 'neigh_op_tnl_3')
// (11, 17, 'neigh_op_lft_3')
// (11, 18, 'neigh_op_bnl_3')

reg n244 = 0;
// (9, 17, 'local_g1_3')
// (9, 17, 'lutff_0/in_2')
// (9, 17, 'sp4_h_r_3')
// (10, 17, 'sp4_h_r_14')
// (11, 17, 'sp4_h_r_27')
// (11, 21, 'local_g3_6')
// (11, 21, 'lutff_3/in_2')
// (11, 21, 'sp4_r_v_b_46')
// (11, 22, 'sp4_r_v_b_35')
// (11, 23, 'sp4_r_v_b_22')
// (11, 24, 'sp4_r_v_b_11')
// (12, 14, 'sp4_r_v_b_38')
// (12, 15, 'sp4_r_v_b_27')
// (12, 16, 'sp4_h_r_8')
// (12, 16, 'sp4_r_v_b_14')
// (12, 17, 'sp4_h_r_38')
// (12, 17, 'sp4_r_v_b_3')
// (12, 20, 'sp4_h_r_11')
// (12, 20, 'sp4_v_t_46')
// (12, 21, 'sp4_v_b_46')
// (12, 22, 'sp4_v_b_35')
// (12, 23, 'sp4_v_b_22')
// (12, 24, 'sp4_v_b_11')
// (13, 13, 'sp4_h_r_3')
// (13, 13, 'sp4_v_t_38')
// (13, 14, 'sp4_v_b_38')
// (13, 15, 'sp4_v_b_27')
// (13, 16, 'sp4_h_r_21')
// (13, 16, 'sp4_v_b_14')
// (13, 17, 'sp4_h_l_38')
// (13, 17, 'sp4_v_b_3')
// (13, 20, 'sp4_h_r_22')
// (14, 13, 'sp4_h_r_14')
// (14, 16, 'sp4_h_r_32')
// (14, 20, 'sp4_h_r_35')
// (15, 12, 'neigh_op_tnr_3')
// (15, 12, 'sp4_r_v_b_38')
// (15, 13, 'local_g2_6')
// (15, 13, 'lutff_0/in_0')
// (15, 13, 'lutff_5/in_3')
// (15, 13, 'neigh_op_rgt_3')
// (15, 13, 'sp4_h_r_27')
// (15, 13, 'sp4_r_v_b_27')
// (15, 13, 'sp4_r_v_b_38')
// (15, 14, 'local_g0_3')
// (15, 14, 'lutff_0/in_1')
// (15, 14, 'lutff_2/in_3')
// (15, 14, 'neigh_op_bnr_3')
// (15, 14, 'sp4_r_v_b_14')
// (15, 14, 'sp4_r_v_b_27')
// (15, 15, 'sp4_r_v_b_14')
// (15, 15, 'sp4_r_v_b_3')
// (15, 16, 'local_g2_5')
// (15, 16, 'lutff_1/in_2')
// (15, 16, 'lutff_2/in_1')
// (15, 16, 'lutff_4/in_1')
// (15, 16, 'lutff_5/in_2')
// (15, 16, 'lutff_7/in_0')
// (15, 16, 'sp4_h_r_45')
// (15, 16, 'sp4_r_v_b_3')
// (15, 17, 'sp4_r_v_b_46')
// (15, 18, 'sp4_r_v_b_35')
// (15, 19, 'sp4_r_v_b_22')
// (15, 20, 'sp4_h_r_46')
// (15, 20, 'sp4_r_v_b_11')
// (16, 4, 'sp12_v_t_22')
// (16, 5, 'sp12_v_b_22')
// (16, 6, 'sp12_v_b_21')
// (16, 7, 'sp12_v_b_18')
// (16, 8, 'sp12_v_b_17')
// (16, 9, 'sp12_v_b_14')
// (16, 10, 'sp12_v_b_13')
// (16, 11, 'sp12_v_b_10')
// (16, 11, 'sp4_v_t_38')
// (16, 12, 'local_g0_3')
// (16, 12, 'local_g1_3')
// (16, 12, 'lutff_3/in_3')
// (16, 12, 'lutff_7/in_0')
// (16, 12, 'neigh_op_top_3')
// (16, 12, 'sp12_v_b_9')
// (16, 12, 'sp4_h_r_8')
// (16, 12, 'sp4_v_b_38')
// (16, 12, 'sp4_v_t_38')
// (16, 13, 'local_g1_3')
// (16, 13, 'lutff_0/in_2')
// (16, 13, 'lutff_2/in_2')
// (16, 13, 'lutff_3/out')
// (16, 13, 'lutff_4/in_2')
// (16, 13, 'lutff_5/in_1')
// (16, 13, 'lutff_7/in_3')
// (16, 13, 'sp12_v_b_6')
// (16, 13, 'sp4_h_r_38')
// (16, 13, 'sp4_v_b_27')
// (16, 13, 'sp4_v_b_38')
// (16, 14, 'local_g1_3')
// (16, 14, 'local_g2_3')
// (16, 14, 'lutff_2/in_2')
// (16, 14, 'lutff_4/in_0')
// (16, 14, 'lutff_6/in_1')
// (16, 14, 'lutff_7/in_2')
// (16, 14, 'neigh_op_bot_3')
// (16, 14, 'sp12_v_b_5')
// (16, 14, 'sp4_v_b_14')
// (16, 14, 'sp4_v_b_27')
// (16, 15, 'local_g0_6')
// (16, 15, 'local_g1_6')
// (16, 15, 'lutff_1/in_3')
// (16, 15, 'lutff_2/in_1')
// (16, 15, 'lutff_4/in_1')
// (16, 15, 'lutff_5/in_2')
// (16, 15, 'sp12_v_b_2')
// (16, 15, 'sp4_h_r_3')
// (16, 15, 'sp4_v_b_14')
// (16, 15, 'sp4_v_b_3')
// (16, 16, 'sp12_v_b_1')
// (16, 16, 'sp4_h_l_45')
// (16, 16, 'sp4_v_b_3')
// (16, 16, 'sp4_v_t_46')
// (16, 17, 'sp4_v_b_46')
// (16, 18, 'sp4_v_b_35')
// (16, 19, 'sp4_v_b_22')
// (16, 20, 'local_g0_3')
// (16, 20, 'lutff_1/in_0')
// (16, 20, 'lutff_2/in_1')
// (16, 20, 'lutff_3/in_2')
// (16, 20, 'lutff_7/in_2')
// (16, 20, 'sp4_h_l_46')
// (16, 20, 'sp4_h_r_5')
// (16, 20, 'sp4_v_b_11')
// (17, 12, 'neigh_op_tnl_3')
// (17, 12, 'sp4_h_r_21')
// (17, 13, 'neigh_op_lft_3')
// (17, 13, 'sp4_h_l_38')
// (17, 14, 'neigh_op_bnl_3')
// (17, 15, 'sp4_h_r_14')
// (17, 20, 'sp4_h_r_16')
// (18, 12, 'sp4_h_r_32')
// (18, 15, 'sp4_h_r_27')
// (18, 20, 'sp4_h_r_29')
// (19, 12, 'local_g2_5')
// (19, 12, 'local_g3_5')
// (19, 12, 'lutff_0/in_0')
// (19, 12, 'lutff_1/in_2')
// (19, 12, 'lutff_2/in_2')
// (19, 12, 'lutff_3/in_1')
// (19, 12, 'lutff_5/in_2')
// (19, 12, 'sp4_h_r_45')
// (19, 15, 'sp4_h_r_38')
// (19, 20, 'local_g2_0')
// (19, 20, 'lutff_6/in_0')
// (19, 20, 'lutff_7/in_1')
// (19, 20, 'sp4_h_r_40')
// (20, 12, 'sp4_h_l_45')
// (20, 15, 'local_g0_3')
// (20, 15, 'local_g1_3')
// (20, 15, 'lutff_0/in_1')
// (20, 15, 'lutff_1/in_0')
// (20, 15, 'lutff_2/in_0')
// (20, 15, 'lutff_3/in_2')
// (20, 15, 'lutff_5/in_1')
// (20, 15, 'lutff_6/in_2')
// (20, 15, 'lutff_7/in_0')
// (20, 15, 'sp4_h_l_38')
// (20, 15, 'sp4_h_r_3')
// (20, 20, 'sp4_h_l_40')
// (21, 15, 'sp4_h_r_14')
// (22, 15, 'local_g2_3')
// (22, 15, 'local_g3_3')
// (22, 15, 'lutff_0/in_2')
// (22, 15, 'lutff_1/in_1')
// (22, 15, 'lutff_2/in_1')
// (22, 15, 'lutff_3/in_1')
// (22, 15, 'lutff_4/in_1')
// (22, 15, 'lutff_5/in_1')
// (22, 15, 'lutff_6/in_2')
// (22, 15, 'lutff_7/in_1')
// (22, 15, 'sp4_h_r_27')
// (23, 15, 'sp4_h_r_38')
// (24, 15, 'sp4_h_l_38')

reg n245 = 0;
// (9, 17, 'sp12_h_r_1')
// (10, 17, 'sp12_h_r_2')
// (11, 17, 'sp12_h_r_5')
// (12, 17, 'sp12_h_r_6')
// (13, 17, 'sp12_h_r_9')
// (14, 17, 'sp12_h_r_10')
// (15, 16, 'neigh_op_tnr_3')
// (15, 17, 'neigh_op_rgt_3')
// (15, 17, 'sp12_h_r_13')
// (15, 18, 'neigh_op_bnr_3')
// (16, 16, 'neigh_op_top_3')
// (16, 17, 'lutff_3/out')
// (16, 17, 'sp12_h_r_14')
// (16, 18, 'neigh_op_bot_3')
// (17, 16, 'neigh_op_tnl_3')
// (17, 17, 'neigh_op_lft_3')
// (17, 17, 'sp12_h_r_17')
// (17, 18, 'neigh_op_bnl_3')
// (18, 17, 'sp12_h_r_18')
// (19, 17, 'sp12_h_r_21')
// (20, 17, 'sp12_h_r_22')
// (21, 17, 'sp12_h_l_22')
// (21, 17, 'sp12_v_t_22')
// (21, 18, 'local_g2_6')
// (21, 18, 'lutff_3/in_1')
// (21, 18, 'sp12_v_b_22')
// (21, 19, 'sp12_v_b_21')
// (21, 20, 'sp12_v_b_18')
// (21, 21, 'sp12_v_b_17')
// (21, 22, 'sp12_v_b_14')
// (21, 23, 'sp12_v_b_13')
// (21, 24, 'sp12_v_b_10')
// (21, 25, 'sp12_v_b_9')
// (21, 26, 'sp12_v_b_6')
// (21, 27, 'sp12_v_b_5')
// (21, 28, 'sp12_v_b_2')
// (21, 29, 'sp12_v_b_1')

wire n246;
// (9, 17, 'sp4_h_r_10')
// (10, 17, 'sp4_h_r_23')
// (11, 17, 'local_g3_2')
// (11, 17, 'lutff_3/in_2')
// (11, 17, 'sp4_h_r_34')
// (12, 16, 'neigh_op_tnr_5')
// (12, 17, 'neigh_op_rgt_5')
// (12, 17, 'sp4_h_r_47')
// (12, 18, 'neigh_op_bnr_5')
// (13, 16, 'neigh_op_top_5')
// (13, 17, 'lutff_5/out')
// (13, 17, 'sp4_h_l_47')
// (13, 17, 'sp4_h_r_10')
// (13, 18, 'neigh_op_bot_5')
// (14, 16, 'neigh_op_tnl_5')
// (14, 17, 'neigh_op_lft_5')
// (14, 17, 'sp4_h_r_23')
// (14, 18, 'neigh_op_bnl_5')
// (15, 17, 'sp4_h_r_34')
// (16, 17, 'sp4_h_r_47')
// (17, 17, 'sp4_h_l_47')

reg n247 = 0;
// (9, 18, 'neigh_op_tnr_0')
// (9, 19, 'neigh_op_rgt_0')
// (9, 20, 'neigh_op_bnr_0')
// (10, 18, 'neigh_op_top_0')
// (10, 19, 'lutff_0/out')
// (10, 20, 'neigh_op_bot_0')
// (11, 18, 'neigh_op_tnl_0')
// (11, 19, 'neigh_op_lft_0')
// (11, 20, 'local_g2_0')
// (11, 20, 'lutff_0/in_0')
// (11, 20, 'neigh_op_bnl_0')

reg n248 = 0;
// (9, 18, 'neigh_op_tnr_1')
// (9, 19, 'neigh_op_rgt_1')
// (9, 20, 'neigh_op_bnr_1')
// (10, 18, 'neigh_op_top_1')
// (10, 19, 'lutff_1/out')
// (10, 20, 'neigh_op_bot_1')
// (11, 18, 'neigh_op_tnl_1')
// (11, 19, 'neigh_op_lft_1')
// (11, 20, 'local_g2_1')
// (11, 20, 'lutff_1/in_0')
// (11, 20, 'neigh_op_bnl_1')

reg n249 = 0;
// (9, 18, 'neigh_op_tnr_2')
// (9, 19, 'neigh_op_rgt_2')
// (9, 20, 'neigh_op_bnr_2')
// (10, 18, 'neigh_op_top_2')
// (10, 19, 'lutff_2/out')
// (10, 20, 'neigh_op_bot_2')
// (11, 18, 'neigh_op_tnl_2')
// (11, 19, 'neigh_op_lft_2')
// (11, 20, 'local_g3_2')
// (11, 20, 'lutff_2/in_3')
// (11, 20, 'neigh_op_bnl_2')

reg n250 = 0;
// (9, 18, 'neigh_op_tnr_3')
// (9, 19, 'neigh_op_rgt_3')
// (9, 20, 'neigh_op_bnr_3')
// (10, 18, 'neigh_op_top_3')
// (10, 19, 'lutff_3/out')
// (10, 20, 'neigh_op_bot_3')
// (11, 18, 'neigh_op_tnl_3')
// (11, 19, 'neigh_op_lft_3')
// (11, 20, 'local_g3_3')
// (11, 20, 'lutff_3/in_3')
// (11, 20, 'neigh_op_bnl_3')

reg n251 = 0;
// (9, 18, 'neigh_op_tnr_4')
// (9, 19, 'neigh_op_rgt_4')
// (9, 20, 'neigh_op_bnr_4')
// (10, 18, 'neigh_op_top_4')
// (10, 19, 'lutff_4/out')
// (10, 20, 'neigh_op_bot_4')
// (11, 18, 'neigh_op_tnl_4')
// (11, 19, 'neigh_op_lft_4')
// (11, 20, 'local_g2_4')
// (11, 20, 'lutff_4/in_0')
// (11, 20, 'neigh_op_bnl_4')

reg n252 = 0;
// (9, 18, 'neigh_op_tnr_5')
// (9, 19, 'neigh_op_rgt_5')
// (9, 20, 'neigh_op_bnr_5')
// (10, 18, 'neigh_op_top_5')
// (10, 19, 'lutff_5/out')
// (10, 20, 'neigh_op_bot_5')
// (11, 18, 'neigh_op_tnl_5')
// (11, 19, 'neigh_op_lft_5')
// (11, 20, 'local_g3_5')
// (11, 20, 'lutff_5/in_3')
// (11, 20, 'neigh_op_bnl_5')

reg n253 = 0;
// (9, 18, 'neigh_op_tnr_6')
// (9, 19, 'neigh_op_rgt_6')
// (9, 20, 'neigh_op_bnr_6')
// (10, 18, 'neigh_op_top_6')
// (10, 19, 'lutff_6/out')
// (10, 20, 'neigh_op_bot_6')
// (11, 18, 'neigh_op_tnl_6')
// (11, 19, 'neigh_op_lft_6')
// (11, 20, 'local_g3_6')
// (11, 20, 'lutff_6/in_3')
// (11, 20, 'neigh_op_bnl_6')

reg n254 = 0;
// (9, 18, 'neigh_op_tnr_7')
// (9, 19, 'neigh_op_rgt_7')
// (9, 20, 'neigh_op_bnr_7')
// (10, 18, 'neigh_op_top_7')
// (10, 19, 'lutff_7/out')
// (10, 20, 'neigh_op_bot_7')
// (11, 18, 'neigh_op_tnl_7')
// (11, 19, 'neigh_op_lft_7')
// (11, 20, 'local_g3_7')
// (11, 20, 'lutff_7/in_3')
// (11, 20, 'neigh_op_bnl_7')

wire n255;
// (9, 18, 'sp12_h_r_0')
// (10, 18, 'sp12_h_r_3')
// (11, 18, 'sp12_h_r_4')
// (12, 17, 'neigh_op_tnr_0')
// (12, 18, 'neigh_op_rgt_0')
// (12, 18, 'sp12_h_r_7')
// (12, 19, 'neigh_op_bnr_0')
// (13, 17, 'neigh_op_top_0')
// (13, 18, 'local_g0_0')
// (13, 18, 'lutff_0/in_2')
// (13, 18, 'lutff_0/out')
// (13, 18, 'sp12_h_r_8')
// (13, 19, 'neigh_op_bot_0')
// (14, 17, 'neigh_op_tnl_0')
// (14, 18, 'neigh_op_lft_0')
// (14, 18, 'sp12_h_r_11')
// (14, 19, 'neigh_op_bnl_0')
// (15, 18, 'sp12_h_r_12')
// (16, 18, 'sp12_h_r_15')
// (17, 18, 'local_g1_0')
// (17, 18, 'lutff_0/in_1')
// (17, 18, 'sp12_h_r_16')
// (18, 18, 'sp12_h_r_19')
// (19, 18, 'sp12_h_r_20')
// (20, 18, 'sp12_h_r_23')
// (21, 18, 'sp12_h_l_23')

reg n256 = 0;
// (9, 18, 'sp12_h_r_1')
// (9, 18, 'sp4_h_r_7')
// (10, 18, 'sp12_h_r_2')
// (10, 18, 'sp4_h_r_18')
// (11, 18, 'local_g0_5')
// (11, 18, 'lutff_1/in_2')
// (11, 18, 'sp12_h_r_5')
// (11, 18, 'sp4_h_r_31')
// (12, 18, 'sp12_h_r_6')
// (12, 18, 'sp4_h_r_42')
// (12, 19, 'sp4_r_v_b_36')
// (12, 19, 'sp4_r_v_b_37')
// (12, 20, 'sp4_r_v_b_24')
// (12, 20, 'sp4_r_v_b_25')
// (12, 21, 'local_g2_5')
// (12, 21, 'lutff_1/in_2')
// (12, 21, 'sp4_r_v_b_12')
// (12, 21, 'sp4_r_v_b_13')
// (12, 22, 'sp4_r_v_b_0')
// (12, 22, 'sp4_r_v_b_1')
// (13, 17, 'local_g2_1')
// (13, 17, 'lutff_6/in_3')
// (13, 17, 'lutff_7/in_0')
// (13, 17, 'neigh_op_tnr_1')
// (13, 18, 'local_g3_1')
// (13, 18, 'lutff_1/in_3')
// (13, 18, 'neigh_op_rgt_1')
// (13, 18, 'sp12_h_r_9')
// (13, 18, 'sp4_h_l_42')
// (13, 18, 'sp4_h_r_7')
// (13, 18, 'sp4_v_t_36')
// (13, 18, 'sp4_v_t_37')
// (13, 19, 'neigh_op_bnr_1')
// (13, 19, 'sp4_v_b_36')
// (13, 19, 'sp4_v_b_37')
// (13, 20, 'sp4_v_b_24')
// (13, 20, 'sp4_v_b_25')
// (13, 21, 'sp4_v_b_12')
// (13, 21, 'sp4_v_b_13')
// (13, 22, 'local_g0_1')
// (13, 22, 'lutff_1/in_2')
// (13, 22, 'sp4_v_b_0')
// (13, 22, 'sp4_v_b_1')
// (14, 17, 'neigh_op_top_1')
// (14, 17, 'sp4_r_v_b_46')
// (14, 18, 'local_g0_2')
// (14, 18, 'lutff_1/in_1')
// (14, 18, 'lutff_1/out')
// (14, 18, 'sp12_h_r_10')
// (14, 18, 'sp4_h_r_18')
// (14, 18, 'sp4_r_v_b_35')
// (14, 19, 'neigh_op_bot_1')
// (14, 19, 'sp4_r_v_b_22')
// (14, 20, 'sp4_r_v_b_11')
// (15, 16, 'sp4_v_t_46')
// (15, 17, 'neigh_op_tnl_1')
// (15, 17, 'sp4_v_b_46')
// (15, 18, 'neigh_op_lft_1')
// (15, 18, 'sp12_h_r_13')
// (15, 18, 'sp4_h_r_31')
// (15, 18, 'sp4_v_b_35')
// (15, 19, 'neigh_op_bnl_1')
// (15, 19, 'sp4_v_b_22')
// (15, 20, 'local_g0_3')
// (15, 20, 'lutff_1/in_2')
// (15, 20, 'sp4_v_b_11')
// (16, 18, 'sp12_h_r_14')
// (16, 18, 'sp4_h_r_42')
// (16, 19, 'sp4_r_v_b_37')
// (16, 20, 'sp4_r_v_b_24')
// (16, 21, 'sp4_r_v_b_13')
// (16, 22, 'sp4_r_v_b_0')
// (17, 18, 'sp12_h_r_17')
// (17, 18, 'sp4_h_l_42')
// (17, 18, 'sp4_v_t_37')
// (17, 19, 'sp4_v_b_37')
// (17, 20, 'sp4_v_b_24')
// (17, 21, 'sp4_v_b_13')
// (17, 22, 'local_g1_0')
// (17, 22, 'lutff_1/in_2')
// (17, 22, 'sp4_v_b_0')
// (18, 18, 'sp12_h_r_18')
// (19, 18, 'sp12_h_r_21')
// (20, 18, 'sp12_h_r_22')
// (21, 18, 'sp12_h_l_22')

wire n257;
// (9, 18, 'sp4_r_v_b_45')
// (9, 19, 'local_g0_3')
// (9, 19, 'lutff_2/in_3')
// (9, 19, 'sp4_r_v_b_32')
// (9, 20, 'sp4_r_v_b_21')
// (9, 21, 'sp4_r_v_b_8')
// (10, 17, 'sp4_v_t_45')
// (10, 18, 'sp4_v_b_45')
// (10, 19, 'sp4_v_b_32')
// (10, 20, 'sp4_v_b_21')
// (10, 21, 'sp4_h_r_3')
// (10, 21, 'sp4_v_b_8')
// (11, 21, 'sp4_h_r_14')
// (12, 20, 'neigh_op_tnr_3')
// (12, 21, 'neigh_op_rgt_3')
// (12, 21, 'sp4_h_r_27')
// (12, 22, 'neigh_op_bnr_3')
// (13, 20, 'neigh_op_top_3')
// (13, 21, 'local_g1_3')
// (13, 21, 'lutff_3/out')
// (13, 21, 'lutff_7/in_1')
// (13, 21, 'sp4_h_r_38')
// (13, 22, 'neigh_op_bot_3')
// (14, 20, 'neigh_op_tnl_3')
// (14, 21, 'neigh_op_lft_3')
// (14, 21, 'sp4_h_l_38')
// (14, 22, 'neigh_op_bnl_3')

wire n258;
// (9, 18, 'sp4_r_v_b_47')
// (9, 19, 'local_g2_2')
// (9, 19, 'lutff_2/in_0')
// (9, 19, 'sp4_r_v_b_34')
// (9, 20, 'sp4_r_v_b_23')
// (9, 21, 'sp4_r_v_b_10')
// (10, 17, 'sp4_v_t_47')
// (10, 18, 'sp4_r_v_b_37')
// (10, 18, 'sp4_v_b_47')
// (10, 19, 'sp4_r_v_b_24')
// (10, 19, 'sp4_v_b_34')
// (10, 20, 'neigh_op_tnr_0')
// (10, 20, 'sp4_r_v_b_13')
// (10, 20, 'sp4_v_b_23')
// (10, 21, 'neigh_op_rgt_0')
// (10, 21, 'sp4_h_r_5')
// (10, 21, 'sp4_r_v_b_0')
// (10, 21, 'sp4_v_b_10')
// (10, 22, 'neigh_op_bnr_0')
// (11, 17, 'local_g0_5')
// (11, 17, 'lutff_4/in_3')
// (11, 17, 'sp4_h_r_5')
// (11, 17, 'sp4_v_t_37')
// (11, 18, 'sp4_v_b_37')
// (11, 19, 'sp4_v_b_24')
// (11, 20, 'neigh_op_top_0')
// (11, 20, 'sp4_v_b_13')
// (11, 21, 'lutff_0/out')
// (11, 21, 'sp4_h_r_16')
// (11, 21, 'sp4_v_b_0')
// (11, 22, 'neigh_op_bot_0')
// (12, 17, 'sp4_h_r_16')
// (12, 20, 'neigh_op_tnl_0')
// (12, 21, 'neigh_op_lft_0')
// (12, 21, 'sp4_h_r_29')
// (12, 22, 'neigh_op_bnl_0')
// (13, 17, 'sp4_h_r_29')
// (13, 21, 'local_g2_0')
// (13, 21, 'lutff_7/in_3')
// (13, 21, 'sp4_h_r_40')
// (14, 17, 'sp4_h_r_40')
// (14, 21, 'sp4_h_l_40')
// (15, 17, 'sp4_h_l_40')

reg n259 = 0;
// (9, 19, 'neigh_op_tnr_0')
// (9, 20, 'neigh_op_rgt_0')
// (9, 21, 'neigh_op_bnr_0')
// (10, 19, 'neigh_op_top_0')
// (10, 20, 'lutff_0/out')
// (10, 21, 'neigh_op_bot_0')
// (11, 19, 'local_g2_0')
// (11, 19, 'lutff_2/in_0')
// (11, 19, 'neigh_op_tnl_0')
// (11, 20, 'neigh_op_lft_0')
// (11, 21, 'neigh_op_bnl_0')

reg n260 = 0;
// (9, 19, 'neigh_op_tnr_1')
// (9, 20, 'neigh_op_rgt_1')
// (9, 21, 'neigh_op_bnr_1')
// (10, 19, 'neigh_op_top_1')
// (10, 20, 'lutff_1/out')
// (10, 21, 'neigh_op_bot_1')
// (11, 19, 'local_g2_1')
// (11, 19, 'lutff_3/in_0')
// (11, 19, 'neigh_op_tnl_1')
// (11, 20, 'neigh_op_lft_1')
// (11, 21, 'neigh_op_bnl_1')

reg n261 = 0;
// (9, 19, 'neigh_op_tnr_2')
// (9, 20, 'neigh_op_rgt_2')
// (9, 21, 'neigh_op_bnr_2')
// (10, 19, 'neigh_op_top_2')
// (10, 20, 'lutff_2/out')
// (10, 21, 'neigh_op_bot_2')
// (11, 19, 'local_g3_2')
// (11, 19, 'lutff_4/in_3')
// (11, 19, 'neigh_op_tnl_2')
// (11, 20, 'neigh_op_lft_2')
// (11, 21, 'neigh_op_bnl_2')

reg n262 = 0;
// (9, 19, 'neigh_op_tnr_3')
// (9, 20, 'neigh_op_rgt_3')
// (9, 21, 'neigh_op_bnr_3')
// (10, 19, 'neigh_op_top_3')
// (10, 20, 'lutff_3/out')
// (10, 21, 'neigh_op_bot_3')
// (11, 19, 'local_g3_3')
// (11, 19, 'lutff_5/in_3')
// (11, 19, 'neigh_op_tnl_3')
// (11, 20, 'neigh_op_lft_3')
// (11, 21, 'neigh_op_bnl_3')

reg n263 = 0;
// (9, 19, 'neigh_op_tnr_4')
// (9, 20, 'neigh_op_rgt_4')
// (9, 21, 'neigh_op_bnr_4')
// (10, 19, 'neigh_op_top_4')
// (10, 20, 'lutff_4/out')
// (10, 21, 'neigh_op_bot_4')
// (11, 19, 'local_g2_4')
// (11, 19, 'lutff_6/in_0')
// (11, 19, 'neigh_op_tnl_4')
// (11, 20, 'neigh_op_lft_4')
// (11, 21, 'neigh_op_bnl_4')

reg n264 = 0;
// (9, 19, 'neigh_op_tnr_5')
// (9, 20, 'neigh_op_rgt_5')
// (9, 21, 'neigh_op_bnr_5')
// (10, 19, 'neigh_op_top_5')
// (10, 20, 'lutff_5/out')
// (10, 21, 'neigh_op_bot_5')
// (11, 19, 'local_g3_5')
// (11, 19, 'lutff_7/in_3')
// (11, 19, 'neigh_op_tnl_5')
// (11, 20, 'neigh_op_lft_5')
// (11, 21, 'neigh_op_bnl_5')

reg n265 = 0;
// (9, 19, 'neigh_op_tnr_6')
// (9, 20, 'neigh_op_rgt_6')
// (9, 21, 'neigh_op_bnr_6')
// (10, 19, 'neigh_op_top_6')
// (10, 20, 'lutff_6/out')
// (10, 21, 'neigh_op_bot_6')
// (11, 19, 'local_g3_6')
// (11, 19, 'lutff_0/in_3')
// (11, 19, 'neigh_op_tnl_6')
// (11, 20, 'neigh_op_lft_6')
// (11, 21, 'neigh_op_bnl_6')

reg n266 = 0;
// (9, 19, 'neigh_op_tnr_7')
// (9, 20, 'neigh_op_rgt_7')
// (9, 21, 'neigh_op_bnr_7')
// (10, 19, 'neigh_op_top_7')
// (10, 20, 'lutff_7/out')
// (10, 21, 'neigh_op_bot_7')
// (11, 19, 'local_g3_7')
// (11, 19, 'lutff_1/in_3')
// (11, 19, 'neigh_op_tnl_7')
// (11, 20, 'neigh_op_lft_7')
// (11, 21, 'neigh_op_bnl_7')

wire n267;
// (9, 19, 'sp12_h_r_0')
// (10, 19, 'sp12_h_r_3')
// (11, 19, 'sp12_h_r_4')
// (12, 18, 'neigh_op_tnr_0')
// (12, 19, 'neigh_op_rgt_0')
// (12, 19, 'sp12_h_r_7')
// (12, 20, 'neigh_op_bnr_0')
// (13, 18, 'neigh_op_top_0')
// (13, 19, 'local_g0_0')
// (13, 19, 'lutff_0/in_2')
// (13, 19, 'lutff_0/out')
// (13, 19, 'sp12_h_r_8')
// (13, 20, 'neigh_op_bot_0')
// (14, 18, 'neigh_op_tnl_0')
// (14, 19, 'neigh_op_lft_0')
// (14, 19, 'sp12_h_r_11')
// (14, 20, 'neigh_op_bnl_0')
// (15, 19, 'sp12_h_r_12')
// (16, 19, 'sp12_h_r_15')
// (17, 19, 'local_g1_0')
// (17, 19, 'lutff_0/in_1')
// (17, 19, 'sp12_h_r_16')
// (18, 19, 'sp12_h_r_19')
// (19, 19, 'sp12_h_r_20')
// (20, 19, 'sp12_h_r_23')
// (21, 19, 'sp12_h_l_23')

reg n268 = 0;
// (9, 19, 'sp12_h_r_1')
// (10, 19, 'sp12_h_r_2')
// (11, 19, 'local_g0_5')
// (11, 19, 'lutff_1/in_2')
// (11, 19, 'sp12_h_r_5')
// (12, 19, 'sp12_h_r_6')
// (12, 20, 'sp4_r_v_b_36')
// (12, 21, 'sp4_r_v_b_25')
// (12, 22, 'local_g2_4')
// (12, 22, 'lutff_1/in_1')
// (12, 22, 'sp4_r_v_b_12')
// (12, 23, 'sp4_r_v_b_1')
// (13, 16, 'sp4_r_v_b_39')
// (13, 17, 'local_g1_2')
// (13, 17, 'lutff_2/in_1')
// (13, 17, 'sp4_r_v_b_26')
// (13, 18, 'neigh_op_tnr_1')
// (13, 18, 'sp4_r_v_b_15')
// (13, 19, 'local_g3_1')
// (13, 19, 'lutff_1/in_3')
// (13, 19, 'neigh_op_rgt_1')
// (13, 19, 'sp12_h_r_9')
// (13, 19, 'sp4_h_r_7')
// (13, 19, 'sp4_r_v_b_2')
// (13, 19, 'sp4_v_t_36')
// (13, 20, 'neigh_op_bnr_1')
// (13, 20, 'sp4_v_b_36')
// (13, 21, 'sp4_v_b_25')
// (13, 22, 'sp4_v_b_12')
// (13, 23, 'local_g1_1')
// (13, 23, 'lutff_1/in_1')
// (13, 23, 'sp4_v_b_1')
// (14, 15, 'sp4_v_t_39')
// (14, 16, 'sp4_v_b_39')
// (14, 17, 'sp4_v_b_26')
// (14, 18, 'neigh_op_top_1')
// (14, 18, 'sp4_r_v_b_46')
// (14, 18, 'sp4_v_b_15')
// (14, 19, 'local_g3_1')
// (14, 19, 'lutff_1/in_1')
// (14, 19, 'lutff_1/out')
// (14, 19, 'sp12_h_r_10')
// (14, 19, 'sp4_h_r_18')
// (14, 19, 'sp4_r_v_b_35')
// (14, 19, 'sp4_v_b_2')
// (14, 20, 'neigh_op_bot_1')
// (14, 20, 'sp4_r_v_b_22')
// (14, 21, 'sp4_r_v_b_11')
// (15, 17, 'sp4_v_t_46')
// (15, 18, 'neigh_op_tnl_1')
// (15, 18, 'sp4_v_b_46')
// (15, 19, 'neigh_op_lft_1')
// (15, 19, 'sp12_h_r_13')
// (15, 19, 'sp4_h_r_31')
// (15, 19, 'sp4_v_b_35')
// (15, 20, 'neigh_op_bnl_1')
// (15, 20, 'sp4_v_b_22')
// (15, 21, 'local_g0_3')
// (15, 21, 'lutff_1/in_2')
// (15, 21, 'sp4_v_b_11')
// (16, 19, 'sp12_h_r_14')
// (16, 19, 'sp4_h_r_42')
// (16, 20, 'sp4_r_v_b_37')
// (16, 21, 'sp4_r_v_b_24')
// (16, 22, 'sp4_r_v_b_13')
// (16, 23, 'sp4_r_v_b_0')
// (17, 19, 'sp12_h_r_17')
// (17, 19, 'sp4_h_l_42')
// (17, 19, 'sp4_v_t_37')
// (17, 20, 'sp4_v_b_37')
// (17, 21, 'sp4_v_b_24')
// (17, 22, 'sp4_v_b_13')
// (17, 23, 'local_g0_0')
// (17, 23, 'lutff_1/in_1')
// (17, 23, 'sp4_v_b_0')
// (18, 19, 'sp12_h_r_18')
// (19, 19, 'sp12_h_r_21')
// (20, 19, 'sp12_h_r_22')
// (21, 19, 'sp12_h_l_22')

reg n269 = 0;
// (9, 19, 'sp4_h_r_5')
// (10, 19, 'sp4_h_r_16')
// (10, 19, 'sp4_h_r_3')
// (11, 19, 'local_g0_6')
// (11, 19, 'lutff_0/in_2')
// (11, 19, 'sp4_h_r_14')
// (11, 19, 'sp4_h_r_29')
// (12, 19, 'sp4_h_r_27')
// (12, 19, 'sp4_h_r_40')
// (12, 20, 'sp4_r_v_b_47')
// (12, 21, 'sp4_r_v_b_34')
// (12, 22, 'local_g3_7')
// (12, 22, 'lutff_0/in_2')
// (12, 22, 'sp4_r_v_b_23')
// (12, 23, 'sp4_r_v_b_10')
// (13, 17, 'local_g3_0')
// (13, 17, 'lutff_2/in_3')
// (13, 17, 'sp4_r_v_b_40')
// (13, 18, 'neigh_op_tnr_0')
// (13, 18, 'sp4_r_v_b_29')
// (13, 19, 'local_g3_0')
// (13, 19, 'lutff_0/in_3')
// (13, 19, 'neigh_op_rgt_0')
// (13, 19, 'sp4_h_l_40')
// (13, 19, 'sp4_h_r_38')
// (13, 19, 'sp4_h_r_5')
// (13, 19, 'sp4_r_v_b_16')
// (13, 19, 'sp4_v_t_47')
// (13, 20, 'neigh_op_bnr_0')
// (13, 20, 'sp4_r_v_b_5')
// (13, 20, 'sp4_v_b_47')
// (13, 21, 'sp4_v_b_34')
// (13, 22, 'sp4_v_b_23')
// (13, 23, 'local_g0_2')
// (13, 23, 'lutff_0/in_2')
// (13, 23, 'sp4_v_b_10')
// (14, 16, 'sp4_v_t_40')
// (14, 17, 'sp4_v_b_40')
// (14, 18, 'neigh_op_top_0')
// (14, 18, 'sp4_r_v_b_44')
// (14, 18, 'sp4_v_b_29')
// (14, 19, 'local_g3_0')
// (14, 19, 'lutff_0/in_1')
// (14, 19, 'lutff_0/out')
// (14, 19, 'sp4_h_l_38')
// (14, 19, 'sp4_h_r_0')
// (14, 19, 'sp4_h_r_16')
// (14, 19, 'sp4_r_v_b_33')
// (14, 19, 'sp4_v_b_16')
// (14, 20, 'neigh_op_bot_0')
// (14, 20, 'sp4_r_v_b_20')
// (14, 20, 'sp4_v_b_5')
// (14, 21, 'sp4_r_v_b_9')
// (15, 17, 'sp4_v_t_44')
// (15, 18, 'neigh_op_tnl_0')
// (15, 18, 'sp4_v_b_44')
// (15, 19, 'neigh_op_lft_0')
// (15, 19, 'sp4_h_r_13')
// (15, 19, 'sp4_h_r_29')
// (15, 19, 'sp4_v_b_33')
// (15, 20, 'neigh_op_bnl_0')
// (15, 20, 'sp4_v_b_20')
// (15, 21, 'local_g1_1')
// (15, 21, 'lutff_0/in_2')
// (15, 21, 'sp4_v_b_9')
// (16, 19, 'sp4_h_r_24')
// (16, 19, 'sp4_h_r_40')
// (17, 19, 'sp4_h_l_40')
// (17, 19, 'sp4_h_r_37')
// (17, 20, 'sp4_r_v_b_37')
// (17, 21, 'sp4_r_v_b_24')
// (17, 22, 'sp4_r_v_b_13')
// (17, 23, 'local_g1_0')
// (17, 23, 'lutff_0/in_1')
// (17, 23, 'sp4_r_v_b_0')
// (18, 19, 'sp4_h_l_37')
// (18, 19, 'sp4_v_t_37')
// (18, 20, 'sp4_v_b_37')
// (18, 21, 'sp4_v_b_24')
// (18, 22, 'sp4_v_b_13')
// (18, 23, 'sp4_v_b_0')

wire n270;
// (9, 20, 'sp12_h_r_1')
// (10, 20, 'sp12_h_r_2')
// (11, 20, 'sp12_h_r_5')
// (12, 20, 'sp12_h_r_6')
// (13, 20, 'sp12_h_r_9')
// (14, 20, 'sp12_h_r_10')
// (15, 19, 'neigh_op_tnr_3')
// (15, 20, 'neigh_op_rgt_3')
// (15, 20, 'sp12_h_r_13')
// (15, 21, 'neigh_op_bnr_3')
// (16, 19, 'neigh_op_top_3')
// (16, 20, 'lutff_3/out')
// (16, 20, 'sp12_h_r_14')
// (16, 21, 'neigh_op_bot_3')
// (17, 19, 'neigh_op_tnl_3')
// (17, 20, 'neigh_op_lft_3')
// (17, 20, 'sp12_h_r_17')
// (17, 21, 'neigh_op_bnl_3')
// (18, 20, 'sp12_h_r_18')
// (19, 20, 'sp12_h_r_21')
// (19, 20, 'sp4_h_r_10')
// (20, 20, 'sp12_h_r_22')
// (20, 20, 'sp4_h_r_23')
// (21, 20, 'local_g2_2')
// (21, 20, 'lutff_global/cen')
// (21, 20, 'sp12_h_l_22')
// (21, 20, 'sp4_h_r_34')
// (22, 20, 'sp4_h_r_47')
// (23, 20, 'sp4_h_l_47')

reg n271 = 0;
// (9, 22, 'neigh_op_tnr_6')
// (9, 23, 'neigh_op_rgt_6')
// (9, 23, 'sp4_h_r_1')
// (9, 24, 'neigh_op_bnr_6')
// (10, 22, 'neigh_op_top_6')
// (10, 23, 'lutff_6/out')
// (10, 23, 'sp4_h_r_12')
// (10, 24, 'neigh_op_bot_6')
// (11, 22, 'neigh_op_tnl_6')
// (11, 23, 'neigh_op_lft_6')
// (11, 23, 'sp4_h_r_25')
// (11, 24, 'neigh_op_bnl_6')
// (12, 20, 'sp4_r_v_b_42')
// (12, 21, 'sp4_r_v_b_31')
// (12, 22, 'sp4_r_v_b_18')
// (12, 23, 'sp4_h_r_36')
// (12, 23, 'sp4_r_v_b_7')
// (13, 19, 'sp4_v_t_42')
// (13, 20, 'sp4_v_b_42')
// (13, 21, 'sp4_v_b_31')
// (13, 22, 'local_g0_2')
// (13, 22, 'lutff_7/in_3')
// (13, 22, 'sp4_v_b_18')
// (13, 23, 'sp4_h_l_36')
// (13, 23, 'sp4_v_b_7')

wire n272;
// (9, 22, 'sp12_h_r_1')
// (10, 22, 'sp12_h_r_2')
// (11, 22, 'sp12_h_r_5')
// (12, 22, 'sp12_h_r_6')
// (13, 22, 'sp12_h_r_9')
// (14, 22, 'sp12_h_r_10')
// (15, 22, 'sp12_h_r_13')
// (16, 22, 'local_g1_6')
// (16, 22, 'lutff_3/in_0')
// (16, 22, 'lutff_4/in_3')
// (16, 22, 'sp12_h_r_14')
// (17, 22, 'sp12_h_r_17')
// (18, 22, 'local_g0_6')
// (18, 22, 'lutff_0/in_0')
// (18, 22, 'lutff_3/in_3')
// (18, 22, 'lutff_5/in_3')
// (18, 22, 'lutff_6/in_0')
// (18, 22, 'lutff_7/in_3')
// (18, 22, 'sp12_h_r_18')
// (18, 22, 'sp4_h_r_6')
// (19, 20, 'local_g2_6')
// (19, 20, 'lutff_0/in_0')
// (19, 20, 'lutff_1/in_3')
// (19, 20, 'lutff_2/in_0')
// (19, 20, 'lutff_3/in_3')
// (19, 20, 'lutff_4/in_0')
// (19, 20, 'sp4_r_v_b_38')
// (19, 21, 'neigh_op_tnr_7')
// (19, 21, 'sp4_r_v_b_27')
// (19, 22, 'neigh_op_rgt_7')
// (19, 22, 'sp12_h_r_21')
// (19, 22, 'sp4_h_r_19')
// (19, 22, 'sp4_r_v_b_14')
// (19, 23, 'local_g0_7')
// (19, 23, 'local_g1_7')
// (19, 23, 'lutff_0/in_1')
// (19, 23, 'lutff_1/in_3')
// (19, 23, 'lutff_2/in_1')
// (19, 23, 'lutff_3/in_3')
// (19, 23, 'lutff_4/in_1')
// (19, 23, 'lutff_5/in_3')
// (19, 23, 'lutff_6/in_1')
// (19, 23, 'lutff_7/in_3')
// (19, 23, 'neigh_op_bnr_7')
// (19, 23, 'sp4_r_v_b_3')
// (20, 19, 'sp4_v_t_38')
// (20, 20, 'sp4_v_b_38')
// (20, 21, 'neigh_op_top_7')
// (20, 21, 'sp4_v_b_27')
// (20, 22, 'lutff_7/out')
// (20, 22, 'sp12_h_r_22')
// (20, 22, 'sp4_h_r_30')
// (20, 22, 'sp4_v_b_14')
// (20, 23, 'neigh_op_bot_7')
// (20, 23, 'sp4_v_b_3')
// (21, 21, 'neigh_op_tnl_7')
// (21, 22, 'neigh_op_lft_7')
// (21, 22, 'sp12_h_l_22')
// (21, 22, 'sp4_h_r_43')
// (21, 23, 'neigh_op_bnl_7')
// (22, 22, 'sp4_h_l_43')

wire n273;
// (9, 22, 'sp4_r_v_b_46')
// (9, 23, 'sp4_r_v_b_35')
// (9, 24, 'sp4_r_v_b_22')
// (9, 25, 'sp4_r_v_b_11')
// (10, 20, 'neigh_op_tnr_3')
// (10, 21, 'neigh_op_rgt_3')
// (10, 21, 'sp4_h_r_11')
// (10, 21, 'sp4_v_t_46')
// (10, 22, 'neigh_op_bnr_3')
// (10, 22, 'sp4_v_b_46')
// (10, 23, 'local_g3_3')
// (10, 23, 'lutff_global/cen')
// (10, 23, 'sp4_v_b_35')
// (10, 24, 'sp4_v_b_22')
// (10, 25, 'sp4_v_b_11')
// (11, 20, 'neigh_op_top_3')
// (11, 21, 'lutff_3/out')
// (11, 21, 'sp4_h_r_22')
// (11, 22, 'local_g1_3')
// (11, 22, 'lutff_global/cen')
// (11, 22, 'neigh_op_bot_3')
// (12, 20, 'neigh_op_tnl_3')
// (12, 21, 'neigh_op_lft_3')
// (12, 21, 'sp4_h_r_35')
// (12, 22, 'neigh_op_bnl_3')
// (13, 21, 'sp4_h_r_46')
// (14, 21, 'sp4_h_l_46')

reg n274 = 0;
// (9, 24, 'sp12_h_r_1')
// (10, 24, 'sp12_h_r_2')
// (11, 24, 'sp12_h_r_5')
// (12, 24, 'sp12_h_r_6')
// (13, 24, 'sp12_h_r_9')
// (14, 24, 'sp12_h_r_10')
// (15, 23, 'neigh_op_tnr_3')
// (15, 24, 'neigh_op_rgt_3')
// (15, 24, 'sp12_h_r_13')
// (15, 25, 'neigh_op_bnr_3')
// (16, 23, 'neigh_op_top_3')
// (16, 24, 'lutff_3/out')
// (16, 24, 'sp12_h_r_14')
// (16, 25, 'neigh_op_bot_3')
// (17, 23, 'neigh_op_tnl_3')
// (17, 24, 'neigh_op_lft_3')
// (17, 24, 'sp12_h_r_17')
// (17, 25, 'neigh_op_bnl_3')
// (18, 24, 'sp12_h_r_18')
// (19, 24, 'sp12_h_r_21')
// (20, 24, 'sp12_h_r_22')
// (21, 24, 'sp12_h_l_22')
// (21, 24, 'sp12_h_r_1')
// (22, 24, 'sp12_h_r_2')
// (23, 24, 'sp12_h_r_5')
// (24, 24, 'sp12_h_r_6')
// (25, 24, 'sp12_h_r_9')
// (26, 24, 'sp12_h_r_10')
// (27, 24, 'sp12_h_r_13')
// (27, 24, 'sp4_h_r_6')
// (28, 24, 'sp12_h_r_14')
// (28, 24, 'sp4_h_r_19')
// (29, 24, 'sp12_h_r_17')
// (29, 24, 'sp4_h_r_30')
// (30, 24, 'sp12_h_r_18')
// (30, 24, 'sp4_h_r_43')
// (30, 25, 'sp4_r_v_b_43')
// (30, 26, 'sp4_r_v_b_30')
// (30, 27, 'sp4_r_v_b_19')
// (30, 28, 'sp4_r_v_b_6')
// (30, 29, 'sp4_r_v_b_43')
// (30, 30, 'sp4_r_v_b_30')
// (30, 31, 'sp4_r_v_b_19')
// (30, 32, 'sp4_r_v_b_6')
// (31, 24, 'sp12_h_r_21')
// (31, 24, 'sp4_h_l_43')
// (31, 24, 'sp4_v_t_43')
// (31, 25, 'sp4_v_b_43')
// (31, 26, 'sp4_v_b_30')
// (31, 27, 'sp4_v_b_19')
// (31, 28, 'sp4_v_b_6')
// (31, 28, 'sp4_v_t_43')
// (31, 29, 'sp4_v_b_43')
// (31, 30, 'sp4_v_b_30')
// (31, 31, 'sp4_v_b_19')
// (31, 32, 'sp4_v_b_6')
// (31, 32, 'sp4_v_t_43')
// (31, 33, 'io_0/D_OUT_0')
// (31, 33, 'local_g1_3')
// (31, 33, 'span4_vert_43')
// (32, 24, 'sp12_h_r_22')
// (33, 24, 'span12_horz_22')

wire io_33_1_1;
// (10, 7, 'sp4_h_r_2')
// (10, 13, 'sp12_h_r_0')
// (11, 7, 'sp4_h_r_15')
// (11, 13, 'sp12_h_r_3')
// (11, 13, 'sp4_h_r_3')
// (12, 7, 'sp4_h_r_26')
// (12, 13, 'sp12_h_r_4')
// (12, 13, 'sp4_h_r_14')
// (13, 7, 'local_g3_7')
// (13, 7, 'lutff_3/in_3')
// (13, 7, 'sp4_h_r_39')
// (13, 8, 'sp4_r_v_b_46')
// (13, 9, 'sp4_r_v_b_35')
// (13, 10, 'sp4_r_v_b_22')
// (13, 11, 'local_g2_3')
// (13, 11, 'lutff_1/in_0')
// (13, 11, 'lutff_2/in_1')
// (13, 11, 'lutff_3/in_2')
// (13, 11, 'lutff_5/in_0')
// (13, 11, 'lutff_6/in_3')
// (13, 11, 'sp4_r_v_b_11')
// (13, 13, 'sp12_h_r_7')
// (13, 13, 'sp4_h_r_27')
// (14, 1, 'sp12_h_r_0')
// (14, 1, 'sp12_v_t_23')
// (14, 2, 'sp12_v_b_23')
// (14, 3, 'sp12_v_b_20')
// (14, 4, 'sp12_v_b_19')
// (14, 5, 'sp12_v_b_16')
// (14, 6, 'sp12_v_b_15')
// (14, 7, 'sp12_v_b_12')
// (14, 7, 'sp4_h_l_39')
// (14, 7, 'sp4_h_r_11')
// (14, 7, 'sp4_v_t_46')
// (14, 8, 'sp12_v_b_11')
// (14, 8, 'sp4_v_b_46')
// (14, 9, 'sp12_v_b_8')
// (14, 9, 'sp4_v_b_35')
// (14, 10, 'sp12_v_b_7')
// (14, 10, 'sp4_r_v_b_44')
// (14, 10, 'sp4_v_b_22')
// (14, 11, 'sp12_v_b_4')
// (14, 11, 'sp4_r_v_b_33')
// (14, 11, 'sp4_v_b_11')
// (14, 12, 'sp12_v_b_3')
// (14, 12, 'sp4_r_v_b_20')
// (14, 13, 'sp12_h_r_8')
// (14, 13, 'sp12_v_b_0')
// (14, 13, 'sp12_v_t_23')
// (14, 13, 'sp4_h_r_38')
// (14, 13, 'sp4_r_v_b_9')
// (14, 14, 'sp12_v_b_23')
// (14, 14, 'sp4_r_v_b_40')
// (14, 15, 'sp12_v_b_20')
// (14, 15, 'sp4_r_v_b_29')
// (14, 16, 'local_g3_0')
// (14, 16, 'local_g3_3')
// (14, 16, 'lutff_5/in_0')
// (14, 16, 'lutff_6/in_2')
// (14, 16, 'sp12_v_b_19')
// (14, 16, 'sp4_r_v_b_16')
// (14, 17, 'sp12_v_b_16')
// (14, 17, 'sp4_r_v_b_5')
// (14, 18, 'sp12_v_b_15')
// (14, 19, 'sp12_v_b_12')
// (14, 20, 'sp12_v_b_11')
// (14, 21, 'sp12_v_b_8')
// (14, 22, 'sp12_v_b_7')
// (14, 23, 'sp12_v_b_4')
// (14, 24, 'sp12_v_b_3')
// (14, 25, 'sp12_v_b_0')
// (15, 1, 'sp12_h_r_3')
// (15, 7, 'local_g0_6')
// (15, 7, 'local_g1_6')
// (15, 7, 'lutff_0/in_0')
// (15, 7, 'lutff_2/in_0')
// (15, 7, 'lutff_6/in_0')
// (15, 7, 'lutff_7/in_0')
// (15, 7, 'sp4_h_r_22')
// (15, 9, 'sp4_v_t_44')
// (15, 10, 'sp4_v_b_44')
// (15, 11, 'sp4_v_b_33')
// (15, 12, 'local_g0_4')
// (15, 12, 'lutff_5/in_1')
// (15, 12, 'sp4_v_b_20')
// (15, 13, 'sp12_h_r_11')
// (15, 13, 'sp4_h_l_38')
// (15, 13, 'sp4_v_b_9')
// (15, 13, 'sp4_v_t_40')
// (15, 14, 'sp4_v_b_40')
// (15, 15, 'sp4_v_b_29')
// (15, 16, 'sp4_v_b_16')
// (15, 17, 'sp4_v_b_5')
// (16, 1, 'sp12_h_r_4')
// (16, 7, 'sp4_h_r_35')
// (16, 13, 'sp12_h_r_12')
// (17, 1, 'sp12_h_r_7')
// (17, 4, 'sp4_r_v_b_43')
// (17, 5, 'sp4_r_v_b_30')
// (17, 6, 'sp4_r_v_b_19')
// (17, 7, 'sp4_h_r_46')
// (17, 7, 'sp4_r_v_b_6')
// (17, 13, 'sp12_h_r_15')
// (18, 1, 'sp12_h_r_0')
// (18, 1, 'sp12_h_r_8')
// (18, 1, 'sp12_v_t_23')
// (18, 2, 'sp12_v_b_23')
// (18, 3, 'sp12_v_b_20')
// (18, 3, 'sp4_v_t_43')
// (18, 4, 'sp12_v_b_19')
// (18, 4, 'sp4_v_b_43')
// (18, 5, 'sp12_v_b_16')
// (18, 5, 'sp4_v_b_30')
// (18, 6, 'sp12_v_b_15')
// (18, 6, 'sp4_v_b_19')
// (18, 7, 'sp12_v_b_12')
// (18, 7, 'sp4_h_l_46')
// (18, 7, 'sp4_v_b_6')
// (18, 8, 'sp12_v_b_11')
// (18, 9, 'sp12_v_b_8')
// (18, 10, 'sp12_v_b_7')
// (18, 11, 'sp12_v_b_4')
// (18, 12, 'sp12_v_b_3')
// (18, 13, 'sp12_h_r_16')
// (18, 13, 'sp12_v_b_0')
// (19, 1, 'sp12_h_r_11')
// (19, 1, 'sp12_h_r_3')
// (19, 13, 'sp12_h_r_19')
// (20, 1, 'sp12_h_r_12')
// (20, 1, 'sp12_h_r_4')
// (20, 13, 'sp12_h_r_20')
// (21, 1, 'sp12_h_r_15')
// (21, 1, 'sp12_h_r_7')
// (21, 13, 'sp12_h_r_23')
// (22, 1, 'sp12_h_r_0')
// (22, 1, 'sp12_h_r_16')
// (22, 1, 'sp12_h_r_8')
// (22, 1, 'sp12_v_t_23')
// (22, 2, 'sp12_v_b_23')
// (22, 3, 'sp12_v_b_20')
// (22, 4, 'sp12_v_b_19')
// (22, 5, 'sp12_v_b_16')
// (22, 6, 'sp12_v_b_15')
// (22, 7, 'sp12_v_b_12')
// (22, 8, 'sp12_v_b_11')
// (22, 9, 'sp12_v_b_8')
// (22, 10, 'sp12_v_b_7')
// (22, 11, 'sp12_v_b_4')
// (22, 12, 'sp12_v_b_3')
// (22, 13, 'sp12_h_l_23')
// (22, 13, 'sp12_v_b_0')
// (23, 1, 'sp12_h_r_11')
// (23, 1, 'sp12_h_r_19')
// (23, 1, 'sp12_h_r_3')
// (24, 1, 'sp12_h_r_12')
// (24, 1, 'sp12_h_r_20')
// (24, 1, 'sp12_h_r_4')
// (25, 1, 'sp12_h_r_15')
// (25, 1, 'sp12_h_r_23')
// (25, 1, 'sp12_h_r_7')
// (26, 1, 'sp12_h_l_23')
// (26, 1, 'sp12_h_r_0')
// (26, 1, 'sp12_h_r_16')
// (26, 1, 'sp12_h_r_8')
// (27, 1, 'sp12_h_r_11')
// (27, 1, 'sp12_h_r_19')
// (27, 1, 'sp12_h_r_3')
// (28, 1, 'sp12_h_r_12')
// (28, 1, 'sp12_h_r_20')
// (28, 1, 'sp12_h_r_4')
// (29, 1, 'sp12_h_r_15')
// (29, 1, 'sp12_h_r_23')
// (29, 1, 'sp12_h_r_7')
// (30, 1, 'sp12_h_l_23')
// (30, 1, 'sp12_h_r_0')
// (30, 1, 'sp12_h_r_16')
// (30, 1, 'sp12_h_r_8')
// (31, 1, 'sp12_h_r_11')
// (31, 1, 'sp12_h_r_19')
// (31, 1, 'sp12_h_r_3')
// (32, 1, 'neigh_op_rgt_2')
// (32, 1, 'neigh_op_rgt_6')
// (32, 1, 'sp12_h_r_12')
// (32, 1, 'sp12_h_r_20')
// (32, 1, 'sp12_h_r_4')
// (32, 2, 'neigh_op_bnr_2')
// (32, 2, 'neigh_op_bnr_6')
// (33, 1, 'io_1/D_IN_0')
// (33, 1, 'io_1/PAD')
// (33, 1, 'span12_horz_12')
// (33, 1, 'span12_horz_20')
// (33, 1, 'span12_horz_4')

wire n276;
// (10, 8, 'neigh_op_tnr_3')
// (10, 9, 'neigh_op_rgt_3')
// (10, 10, 'neigh_op_bnr_3')
// (11, 8, 'neigh_op_top_3')
// (11, 9, 'local_g0_3')
// (11, 9, 'lutff_3/out')
// (11, 9, 'lutff_6/in_1')
// (11, 10, 'neigh_op_bot_3')
// (12, 8, 'neigh_op_tnl_3')
// (12, 9, 'neigh_op_lft_3')
// (12, 10, 'neigh_op_bnl_3')

wire n277;
// (10, 8, 'neigh_op_tnr_4')
// (10, 9, 'local_g3_4')
// (10, 9, 'lutff_0/in_3')
// (10, 9, 'neigh_op_rgt_4')
// (10, 10, 'local_g1_4')
// (10, 10, 'lutff_0/in_1')
// (10, 10, 'neigh_op_bnr_4')
// (11, 8, 'neigh_op_top_4')
// (11, 9, 'lutff_4/out')
// (11, 10, 'neigh_op_bot_4')
// (12, 8, 'neigh_op_tnl_4')
// (12, 9, 'neigh_op_lft_4')
// (12, 10, 'neigh_op_bnl_4')

reg n278 = 0;
// (10, 8, 'neigh_op_tnr_5')
// (10, 9, 'neigh_op_rgt_5')
// (10, 10, 'neigh_op_bnr_5')
// (11, 8, 'neigh_op_top_5')
// (11, 8, 'sp4_r_v_b_38')
// (11, 9, 'local_g2_5')
// (11, 9, 'lutff_5/in_2')
// (11, 9, 'lutff_5/out')
// (11, 9, 'sp4_r_v_b_27')
// (11, 10, 'neigh_op_bot_5')
// (11, 10, 'sp4_r_v_b_14')
// (11, 11, 'sp4_r_v_b_3')
// (12, 7, 'sp4_v_t_38')
// (12, 8, 'neigh_op_tnl_5')
// (12, 8, 'sp4_v_b_38')
// (12, 9, 'neigh_op_lft_5')
// (12, 9, 'sp4_v_b_27')
// (12, 10, 'neigh_op_bnl_5')
// (12, 10, 'sp4_v_b_14')
// (12, 11, 'sp4_h_r_3')
// (12, 11, 'sp4_v_b_3')
// (13, 11, 'sp4_h_r_14')
// (14, 11, 'sp4_h_r_27')
// (15, 11, 'local_g3_6')
// (15, 11, 'lutff_4/in_3')
// (15, 11, 'sp4_h_r_38')
// (16, 11, 'sp4_h_l_38')

wire n279;
// (10, 8, 'neigh_op_tnr_6')
// (10, 9, 'local_g2_6')
// (10, 9, 'local_g3_6')
// (10, 9, 'lutff_0/in_0')
// (10, 9, 'lutff_1/in_0')
// (10, 9, 'lutff_5/in_0')
// (10, 9, 'neigh_op_rgt_6')
// (10, 10, 'neigh_op_bnr_6')
// (11, 8, 'neigh_op_top_6')
// (11, 9, 'local_g2_6')
// (11, 9, 'lutff_5/in_3')
// (11, 9, 'lutff_6/out')
// (11, 10, 'neigh_op_bot_6')
// (12, 8, 'neigh_op_tnl_6')
// (12, 9, 'neigh_op_lft_6')
// (12, 10, 'neigh_op_bnl_6')

reg n280 = 0;
// (10, 8, 'sp4_r_v_b_45')
// (10, 9, 'sp4_r_v_b_32')
// (10, 10, 'neigh_op_tnr_4')
// (10, 10, 'sp4_r_v_b_21')
// (10, 11, 'neigh_op_rgt_4')
// (10, 11, 'sp4_r_v_b_8')
// (10, 12, 'neigh_op_bnr_4')
// (11, 7, 'sp4_v_t_45')
// (11, 8, 'sp4_v_b_45')
// (11, 9, 'local_g2_0')
// (11, 9, 'lutff_1/in_3')
// (11, 9, 'sp4_v_b_32')
// (11, 10, 'local_g1_4')
// (11, 10, 'lutff_2/in_3')
// (11, 10, 'neigh_op_top_4')
// (11, 10, 'sp4_v_b_21')
// (11, 11, 'local_g3_4')
// (11, 11, 'lutff_4/in_1')
// (11, 11, 'lutff_4/out')
// (11, 11, 'sp4_v_b_8')
// (11, 12, 'neigh_op_bot_4')
// (12, 10, 'neigh_op_tnl_4')
// (12, 11, 'neigh_op_lft_4')
// (12, 12, 'neigh_op_bnl_4')

reg n281 = 0;
// (10, 8, 'sp4_r_v_b_47')
// (10, 9, 'sp4_r_v_b_34')
// (10, 10, 'neigh_op_tnr_5')
// (10, 10, 'sp4_r_v_b_23')
// (10, 11, 'neigh_op_rgt_5')
// (10, 11, 'sp4_r_v_b_10')
// (10, 12, 'neigh_op_bnr_5')
// (11, 7, 'sp4_v_t_47')
// (11, 8, 'sp4_v_b_47')
// (11, 9, 'local_g3_2')
// (11, 9, 'lutff_1/in_0')
// (11, 9, 'sp4_v_b_34')
// (11, 10, 'local_g0_5')
// (11, 10, 'lutff_2/in_1')
// (11, 10, 'neigh_op_top_5')
// (11, 10, 'sp4_v_b_23')
// (11, 11, 'local_g1_5')
// (11, 11, 'lutff_5/in_1')
// (11, 11, 'lutff_5/out')
// (11, 11, 'sp4_v_b_10')
// (11, 12, 'neigh_op_bot_5')
// (12, 10, 'neigh_op_tnl_5')
// (12, 11, 'neigh_op_lft_5')
// (12, 12, 'neigh_op_bnl_5')

wire n282;
// (10, 9, 'neigh_op_tnr_0')
// (10, 10, 'neigh_op_rgt_0')
// (10, 11, 'neigh_op_bnr_0')
// (11, 9, 'neigh_op_top_0')
// (11, 10, 'local_g2_0')
// (11, 10, 'lutff_0/out')
// (11, 10, 'lutff_7/in_3')
// (11, 11, 'local_g0_0')
// (11, 11, 'local_g1_0')
// (11, 11, 'lutff_2/in_0')
// (11, 11, 'lutff_3/in_0')
// (11, 11, 'lutff_4/in_0')
// (11, 11, 'lutff_5/in_0')
// (11, 11, 'lutff_6/in_0')
// (11, 11, 'lutff_7/in_0')
// (11, 11, 'neigh_op_bot_0')
// (12, 9, 'neigh_op_tnl_0')
// (12, 10, 'neigh_op_lft_0')
// (12, 11, 'neigh_op_bnl_0')

reg n283 = 0;
// (10, 9, 'neigh_op_tnr_1')
// (10, 10, 'neigh_op_rgt_1')
// (10, 11, 'neigh_op_bnr_1')
// (11, 9, 'neigh_op_top_1')
// (11, 10, 'local_g3_1')
// (11, 10, 'lutff_1/out')
// (11, 10, 'lutff_3/in_3')
// (11, 11, 'local_g1_1')
// (11, 11, 'lutff_1/in_1')
// (11, 11, 'neigh_op_bot_1')
// (12, 9, 'neigh_op_tnl_1')
// (12, 10, 'neigh_op_lft_1')
// (12, 11, 'neigh_op_bnl_1')

wire n284;
// (10, 9, 'neigh_op_tnr_3')
// (10, 10, 'neigh_op_rgt_3')
// (10, 11, 'neigh_op_bnr_3')
// (11, 9, 'neigh_op_top_3')
// (11, 10, 'local_g0_3')
// (11, 10, 'lutff_0/in_3')
// (11, 10, 'lutff_1/in_0')
// (11, 10, 'lutff_3/out')
// (11, 10, 'lutff_7/in_0')
// (11, 11, 'neigh_op_bot_3')
// (12, 9, 'neigh_op_tnl_3')
// (12, 10, 'neigh_op_lft_3')
// (12, 11, 'neigh_op_bnl_3')

reg n285 = 0;
// (10, 9, 'neigh_op_tnr_7')
// (10, 10, 'neigh_op_rgt_7')
// (10, 11, 'neigh_op_bnr_7')
// (11, 9, 'neigh_op_top_7')
// (11, 10, 'lutff_7/out')
// (11, 11, 'local_g0_7')
// (11, 11, 'lutff_0/in_1')
// (11, 11, 'neigh_op_bot_7')
// (12, 9, 'neigh_op_tnl_7')
// (12, 10, 'neigh_op_lft_7')
// (12, 11, 'neigh_op_bnl_7')

reg n286 = 0;
// (10, 9, 'sp4_r_v_b_46')
// (10, 10, 'neigh_op_tnr_3')
// (10, 10, 'sp4_r_v_b_35')
// (10, 11, 'neigh_op_rgt_3')
// (10, 11, 'sp4_r_v_b_22')
// (10, 12, 'neigh_op_bnr_3')
// (10, 12, 'sp4_r_v_b_11')
// (11, 8, 'sp4_v_t_46')
// (11, 9, 'sp4_r_v_b_47')
// (11, 9, 'sp4_v_b_46')
// (11, 10, 'local_g2_3')
// (11, 10, 'lutff_3/in_0')
// (11, 10, 'neigh_op_top_3')
// (11, 10, 'sp4_r_v_b_34')
// (11, 10, 'sp4_v_b_35')
// (11, 11, 'local_g1_3')
// (11, 11, 'lutff_3/in_1')
// (11, 11, 'lutff_3/out')
// (11, 11, 'sp4_r_v_b_23')
// (11, 11, 'sp4_v_b_22')
// (11, 12, 'neigh_op_bot_3')
// (11, 12, 'sp4_r_v_b_10')
// (11, 12, 'sp4_v_b_11')
// (12, 8, 'sp4_v_t_47')
// (12, 9, 'local_g2_7')
// (12, 9, 'lutff_3/in_2')
// (12, 9, 'sp4_v_b_47')
// (12, 10, 'neigh_op_tnl_3')
// (12, 10, 'sp4_v_b_34')
// (12, 11, 'neigh_op_lft_3')
// (12, 11, 'sp4_v_b_23')
// (12, 12, 'neigh_op_bnl_3')
// (12, 12, 'sp4_v_b_10')

wire n287;
// (10, 10, 'lutff_0/cout')
// (10, 10, 'lutff_1/in_3')

wire n288;
// (10, 10, 'lutff_1/cout')
// (10, 10, 'lutff_2/in_3')

wire n289;
// (10, 10, 'lutff_2/cout')
// (10, 10, 'lutff_3/in_3')

wire n290;
// (10, 10, 'lutff_3/cout')
// (10, 10, 'lutff_4/in_3')

wire n291;
// (10, 10, 'lutff_7/cout')
// (10, 11, 'carry_in')
// (10, 11, 'carry_in_mux')
// (10, 11, 'lutff_0/in_3')

wire n292;
// (10, 10, 'neigh_op_tnr_0')
// (10, 11, 'neigh_op_rgt_0')
// (10, 12, 'neigh_op_bnr_0')
// (11, 10, 'local_g1_0')
// (11, 10, 'lutff_7/in_2')
// (11, 10, 'neigh_op_top_0')
// (11, 11, 'lutff_0/out')
// (11, 12, 'neigh_op_bot_0')
// (12, 10, 'neigh_op_tnl_0')
// (12, 11, 'neigh_op_lft_0')
// (12, 12, 'neigh_op_bnl_0')

wire n293;
// (10, 10, 'neigh_op_tnr_1')
// (10, 11, 'neigh_op_rgt_1')
// (10, 12, 'neigh_op_bnr_1')
// (11, 10, 'local_g1_1')
// (11, 10, 'lutff_1/in_3')
// (11, 10, 'neigh_op_top_1')
// (11, 11, 'lutff_1/out')
// (11, 12, 'neigh_op_bot_1')
// (12, 10, 'neigh_op_tnl_1')
// (12, 11, 'neigh_op_lft_1')
// (12, 12, 'neigh_op_bnl_1')

reg n294 = 0;
// (10, 10, 'neigh_op_tnr_2')
// (10, 11, 'neigh_op_rgt_2')
// (10, 12, 'neigh_op_bnr_2')
// (11, 9, 'sp4_r_v_b_45')
// (11, 10, 'local_g0_2')
// (11, 10, 'lutff_3/in_1')
// (11, 10, 'neigh_op_top_2')
// (11, 10, 'sp4_r_v_b_32')
// (11, 11, 'local_g1_2')
// (11, 11, 'lutff_2/in_1')
// (11, 11, 'lutff_2/out')
// (11, 11, 'sp4_r_v_b_21')
// (11, 12, 'neigh_op_bot_2')
// (11, 12, 'sp4_r_v_b_8')
// (12, 8, 'sp4_v_t_45')
// (12, 9, 'local_g2_5')
// (12, 9, 'lutff_3/in_0')
// (12, 9, 'sp4_v_b_45')
// (12, 10, 'neigh_op_tnl_2')
// (12, 10, 'sp4_v_b_32')
// (12, 11, 'neigh_op_lft_2')
// (12, 11, 'sp4_v_b_21')
// (12, 12, 'neigh_op_bnl_2')
// (12, 12, 'sp4_v_b_8')

reg n295 = 0;
// (10, 10, 'neigh_op_tnr_6')
// (10, 11, 'neigh_op_rgt_6')
// (10, 12, 'neigh_op_bnr_6')
// (11, 9, 'sp4_r_v_b_37')
// (11, 10, 'local_g0_6')
// (11, 10, 'lutff_2/in_0')
// (11, 10, 'neigh_op_top_6')
// (11, 10, 'sp4_r_v_b_24')
// (11, 11, 'local_g1_6')
// (11, 11, 'lutff_6/in_1')
// (11, 11, 'lutff_6/out')
// (11, 11, 'sp4_r_v_b_13')
// (11, 12, 'neigh_op_bot_6')
// (11, 12, 'sp4_r_v_b_0')
// (12, 8, 'sp4_v_t_37')
// (12, 9, 'local_g3_5')
// (12, 9, 'lutff_3/in_3')
// (12, 9, 'sp4_v_b_37')
// (12, 10, 'neigh_op_tnl_6')
// (12, 10, 'sp4_v_b_24')
// (12, 11, 'neigh_op_lft_6')
// (12, 11, 'sp4_v_b_13')
// (12, 12, 'neigh_op_bnl_6')
// (12, 12, 'sp4_v_b_0')

reg n296 = 0;
// (10, 10, 'neigh_op_tnr_7')
// (10, 11, 'neigh_op_rgt_7')
// (10, 12, 'neigh_op_bnr_7')
// (11, 9, 'sp4_r_v_b_39')
// (11, 10, 'local_g1_7')
// (11, 10, 'lutff_2/in_2')
// (11, 10, 'neigh_op_top_7')
// (11, 10, 'sp4_r_v_b_26')
// (11, 11, 'local_g1_7')
// (11, 11, 'lutff_7/in_1')
// (11, 11, 'lutff_7/out')
// (11, 11, 'sp4_r_v_b_15')
// (11, 12, 'neigh_op_bot_7')
// (11, 12, 'sp4_r_v_b_2')
// (12, 8, 'sp4_v_t_39')
// (12, 9, 'local_g3_7')
// (12, 9, 'lutff_3/in_1')
// (12, 9, 'sp4_v_b_39')
// (12, 10, 'neigh_op_tnl_7')
// (12, 10, 'sp4_v_b_26')
// (12, 11, 'neigh_op_lft_7')
// (12, 11, 'sp4_v_b_15')
// (12, 12, 'neigh_op_bnl_7')
// (12, 12, 'sp4_v_b_2')

reg n297 = 0;
// (10, 12, 'neigh_op_tnr_0')
// (10, 12, 'sp4_r_v_b_45')
// (10, 13, 'neigh_op_rgt_0')
// (10, 13, 'sp4_r_v_b_32')
// (10, 14, 'neigh_op_bnr_0')
// (10, 14, 'sp4_r_v_b_21')
// (10, 15, 'sp4_r_v_b_8')
// (11, 11, 'sp4_v_t_45')
// (11, 12, 'neigh_op_top_0')
// (11, 12, 'sp4_v_b_45')
// (11, 13, 'lutff_0/out')
// (11, 13, 'sp4_v_b_32')
// (11, 14, 'neigh_op_bot_0')
// (11, 14, 'sp4_v_b_21')
// (11, 15, 'local_g0_0')
// (11, 15, 'lutff_2/in_2')
// (11, 15, 'sp4_v_b_8')
// (12, 12, 'neigh_op_tnl_0')
// (12, 13, 'neigh_op_lft_0')
// (12, 14, 'neigh_op_bnl_0')

reg n298 = 0;
// (10, 12, 'neigh_op_tnr_1')
// (10, 12, 'sp4_r_v_b_47')
// (10, 13, 'neigh_op_rgt_1')
// (10, 13, 'sp4_r_v_b_34')
// (10, 14, 'neigh_op_bnr_1')
// (10, 14, 'sp4_r_v_b_23')
// (10, 15, 'sp4_r_v_b_10')
// (11, 11, 'sp4_v_t_47')
// (11, 12, 'neigh_op_top_1')
// (11, 12, 'sp4_v_b_47')
// (11, 13, 'lutff_1/out')
// (11, 13, 'sp4_v_b_34')
// (11, 14, 'neigh_op_bot_1')
// (11, 14, 'sp4_v_b_23')
// (11, 15, 'local_g1_2')
// (11, 15, 'lutff_3/in_2')
// (11, 15, 'sp4_v_b_10')
// (12, 12, 'neigh_op_tnl_1')
// (12, 13, 'neigh_op_lft_1')
// (12, 14, 'neigh_op_bnl_1')

reg n299 = 0;
// (10, 12, 'neigh_op_tnr_2')
// (10, 13, 'neigh_op_rgt_2')
// (10, 13, 'sp4_r_v_b_36')
// (10, 14, 'neigh_op_bnr_2')
// (10, 14, 'sp4_r_v_b_25')
// (10, 15, 'sp4_r_v_b_12')
// (10, 16, 'sp4_r_v_b_1')
// (11, 12, 'neigh_op_top_2')
// (11, 12, 'sp4_v_t_36')
// (11, 13, 'lutff_2/out')
// (11, 13, 'sp4_v_b_36')
// (11, 14, 'neigh_op_bot_2')
// (11, 14, 'sp4_v_b_25')
// (11, 15, 'local_g0_4')
// (11, 15, 'lutff_4/in_2')
// (11, 15, 'sp4_v_b_12')
// (11, 16, 'sp4_v_b_1')
// (12, 12, 'neigh_op_tnl_2')
// (12, 13, 'neigh_op_lft_2')
// (12, 14, 'neigh_op_bnl_2')

reg n300 = 0;
// (10, 12, 'neigh_op_tnr_3')
// (10, 13, 'neigh_op_rgt_3')
// (10, 14, 'neigh_op_bnr_3')
// (11, 12, 'neigh_op_top_3')
// (11, 13, 'lutff_3/out')
// (11, 13, 'sp4_r_v_b_39')
// (11, 14, 'neigh_op_bot_3')
// (11, 14, 'sp4_r_v_b_26')
// (11, 15, 'local_g2_7')
// (11, 15, 'lutff_5/in_2')
// (11, 15, 'sp4_r_v_b_15')
// (11, 16, 'sp4_r_v_b_2')
// (12, 12, 'neigh_op_tnl_3')
// (12, 12, 'sp4_v_t_39')
// (12, 13, 'neigh_op_lft_3')
// (12, 13, 'sp4_v_b_39')
// (12, 14, 'neigh_op_bnl_3')
// (12, 14, 'sp4_v_b_26')
// (12, 15, 'sp4_v_b_15')
// (12, 16, 'sp4_v_b_2')

reg n301 = 0;
// (10, 12, 'neigh_op_tnr_4')
// (10, 13, 'neigh_op_rgt_4')
// (10, 14, 'neigh_op_bnr_4')
// (11, 12, 'neigh_op_top_4')
// (11, 13, 'lutff_4/out')
// (11, 13, 'sp4_r_v_b_41')
// (11, 14, 'neigh_op_bot_4')
// (11, 14, 'sp4_r_v_b_28')
// (11, 15, 'local_g3_1')
// (11, 15, 'lutff_6/in_2')
// (11, 15, 'sp4_r_v_b_17')
// (11, 16, 'sp4_r_v_b_4')
// (12, 12, 'neigh_op_tnl_4')
// (12, 12, 'sp4_v_t_41')
// (12, 13, 'neigh_op_lft_4')
// (12, 13, 'sp4_v_b_41')
// (12, 14, 'neigh_op_bnl_4')
// (12, 14, 'sp4_v_b_28')
// (12, 15, 'sp4_v_b_17')
// (12, 16, 'sp4_v_b_4')

reg n302 = 0;
// (10, 12, 'neigh_op_tnr_5')
// (10, 13, 'neigh_op_rgt_5')
// (10, 13, 'sp4_r_v_b_42')
// (10, 14, 'neigh_op_bnr_5')
// (10, 14, 'sp4_r_v_b_31')
// (10, 15, 'sp4_r_v_b_18')
// (10, 16, 'sp4_r_v_b_7')
// (11, 12, 'neigh_op_top_5')
// (11, 12, 'sp4_v_t_42')
// (11, 13, 'lutff_5/out')
// (11, 13, 'sp4_v_b_42')
// (11, 14, 'neigh_op_bot_5')
// (11, 14, 'sp4_v_b_31')
// (11, 15, 'local_g0_2')
// (11, 15, 'lutff_7/in_1')
// (11, 15, 'sp4_v_b_18')
// (11, 16, 'sp4_v_b_7')
// (12, 12, 'neigh_op_tnl_5')
// (12, 13, 'neigh_op_lft_5')
// (12, 14, 'neigh_op_bnl_5')

reg n303 = 0;
// (10, 12, 'neigh_op_tnr_6')
// (10, 13, 'neigh_op_rgt_6')
// (10, 14, 'neigh_op_bnr_6')
// (11, 12, 'neigh_op_top_6')
// (11, 13, 'lutff_6/out')
// (11, 13, 'sp4_r_v_b_45')
// (11, 14, 'neigh_op_bot_6')
// (11, 14, 'sp4_r_v_b_32')
// (11, 15, 'local_g3_5')
// (11, 15, 'lutff_0/in_2')
// (11, 15, 'sp4_r_v_b_21')
// (11, 16, 'sp4_r_v_b_8')
// (12, 12, 'neigh_op_tnl_6')
// (12, 12, 'sp4_v_t_45')
// (12, 13, 'neigh_op_lft_6')
// (12, 13, 'sp4_v_b_45')
// (12, 14, 'neigh_op_bnl_6')
// (12, 14, 'sp4_v_b_32')
// (12, 15, 'sp4_v_b_21')
// (12, 16, 'sp4_v_b_8')

reg n304 = 0;
// (10, 12, 'neigh_op_tnr_7')
// (10, 13, 'neigh_op_rgt_7')
// (10, 13, 'sp4_r_v_b_46')
// (10, 14, 'neigh_op_bnr_7')
// (10, 14, 'sp4_r_v_b_35')
// (10, 15, 'sp4_r_v_b_22')
// (10, 16, 'sp4_r_v_b_11')
// (11, 12, 'neigh_op_top_7')
// (11, 12, 'sp4_v_t_46')
// (11, 13, 'lutff_7/out')
// (11, 13, 'sp4_v_b_46')
// (11, 14, 'neigh_op_bot_7')
// (11, 14, 'sp4_v_b_35')
// (11, 15, 'local_g1_6')
// (11, 15, 'lutff_1/in_2')
// (11, 15, 'sp4_v_b_22')
// (11, 16, 'sp4_v_b_11')
// (12, 12, 'neigh_op_tnl_7')
// (12, 13, 'neigh_op_lft_7')
// (12, 14, 'neigh_op_bnl_7')

wire n305;
// (10, 13, 'carry_in_mux')
// (10, 13, 'lutff_0/in_3')

wire n306;
// (10, 13, 'lutff_0/cout')
// (10, 13, 'lutff_1/in_3')

wire n307;
// (10, 13, 'lutff_1/cout')
// (10, 13, 'lutff_2/in_3')

wire n308;
// (10, 13, 'lutff_2/cout')
// (10, 13, 'lutff_3/in_3')

wire n309;
// (10, 13, 'lutff_3/cout')
// (10, 13, 'lutff_4/in_3')

wire n310;
// (10, 13, 'lutff_4/cout')
// (10, 13, 'lutff_5/in_3')

wire n311;
// (10, 13, 'lutff_5/cout')
// (10, 13, 'lutff_6/in_3')

wire n312;
// (10, 13, 'lutff_6/cout')
// (10, 13, 'lutff_7/in_3')

wire n313;
// (10, 13, 'neigh_op_tnr_1')
// (10, 14, 'neigh_op_rgt_1')
// (10, 15, 'neigh_op_bnr_1')
// (11, 13, 'neigh_op_top_1')
// (11, 14, 'lutff_1/out')
// (11, 15, 'neigh_op_bot_1')
// (12, 13, 'neigh_op_tnl_1')
// (12, 14, 'local_g0_1')
// (12, 14, 'lutff_1/in_2')
// (12, 14, 'neigh_op_lft_1')
// (12, 15, 'neigh_op_bnl_1')

wire n314;
// (10, 13, 'neigh_op_tnr_2')
// (10, 14, 'neigh_op_rgt_2')
// (10, 15, 'neigh_op_bnr_2')
// (11, 13, 'neigh_op_top_2')
// (11, 14, 'lutff_2/out')
// (11, 15, 'neigh_op_bot_2')
// (12, 13, 'neigh_op_tnl_2')
// (12, 14, 'local_g0_2')
// (12, 14, 'lutff_2/in_2')
// (12, 14, 'neigh_op_lft_2')
// (12, 15, 'neigh_op_bnl_2')

wire n315;
// (10, 13, 'neigh_op_tnr_3')
// (10, 14, 'neigh_op_rgt_3')
// (10, 15, 'neigh_op_bnr_3')
// (11, 13, 'neigh_op_top_3')
// (11, 14, 'lutff_3/out')
// (11, 15, 'neigh_op_bot_3')
// (12, 13, 'neigh_op_tnl_3')
// (12, 14, 'local_g0_3')
// (12, 14, 'lutff_3/in_2')
// (12, 14, 'neigh_op_lft_3')
// (12, 15, 'neigh_op_bnl_3')

wire n316;
// (10, 13, 'neigh_op_tnr_4')
// (10, 14, 'neigh_op_rgt_4')
// (10, 15, 'neigh_op_bnr_4')
// (11, 13, 'neigh_op_top_4')
// (11, 14, 'lutff_4/out')
// (11, 15, 'neigh_op_bot_4')
// (12, 13, 'neigh_op_tnl_4')
// (12, 14, 'local_g0_4')
// (12, 14, 'lutff_4/in_2')
// (12, 14, 'neigh_op_lft_4')
// (12, 15, 'neigh_op_bnl_4')

wire n317;
// (10, 13, 'neigh_op_tnr_5')
// (10, 14, 'neigh_op_rgt_5')
// (10, 15, 'neigh_op_bnr_5')
// (11, 13, 'neigh_op_top_5')
// (11, 14, 'lutff_5/out')
// (11, 15, 'neigh_op_bot_5')
// (12, 13, 'neigh_op_tnl_5')
// (12, 14, 'local_g0_5')
// (12, 14, 'lutff_5/in_2')
// (12, 14, 'neigh_op_lft_5')
// (12, 15, 'neigh_op_bnl_5')

wire n318;
// (10, 13, 'neigh_op_tnr_6')
// (10, 14, 'neigh_op_rgt_6')
// (10, 15, 'neigh_op_bnr_6')
// (11, 13, 'neigh_op_top_6')
// (11, 14, 'lutff_6/out')
// (11, 15, 'neigh_op_bot_6')
// (12, 13, 'neigh_op_tnl_6')
// (12, 14, 'local_g0_6')
// (12, 14, 'lutff_6/in_2')
// (12, 14, 'neigh_op_lft_6')
// (12, 15, 'neigh_op_bnl_6')

wire n319;
// (10, 13, 'neigh_op_tnr_7')
// (10, 14, 'neigh_op_rgt_7')
// (10, 15, 'neigh_op_bnr_7')
// (11, 13, 'neigh_op_top_7')
// (11, 14, 'lutff_7/out')
// (11, 15, 'neigh_op_bot_7')
// (12, 13, 'neigh_op_tnl_7')
// (12, 14, 'local_g0_7')
// (12, 14, 'lutff_7/in_2')
// (12, 14, 'neigh_op_lft_7')
// (12, 15, 'neigh_op_bnl_7')

wire n320;
// (10, 13, 'sp4_h_r_1')
// (11, 13, 'sp4_h_r_12')
// (12, 12, 'neigh_op_tnr_2')
// (12, 13, 'neigh_op_rgt_2')
// (12, 13, 'sp4_h_r_25')
// (12, 14, 'neigh_op_bnr_2')
// (13, 12, 'neigh_op_top_2')
// (13, 13, 'lutff_2/out')
// (13, 13, 'sp4_h_r_36')
// (13, 14, 'neigh_op_bot_2')
// (13, 14, 'sp4_r_v_b_43')
// (13, 15, 'sp4_r_v_b_30')
// (13, 16, 'sp4_r_v_b_19')
// (13, 17, 'sp4_r_v_b_6')
// (14, 12, 'neigh_op_tnl_2')
// (14, 13, 'neigh_op_lft_2')
// (14, 13, 'sp4_h_l_36')
// (14, 13, 'sp4_v_t_43')
// (14, 14, 'neigh_op_bnl_2')
// (14, 14, 'sp4_v_b_43')
// (14, 15, 'sp4_v_b_30')
// (14, 16, 'local_g0_3')
// (14, 16, 'lutff_6/in_1')
// (14, 16, 'sp4_v_b_19')
// (14, 17, 'sp4_v_b_6')

wire n321;
// (10, 13, 'sp4_h_r_10')
// (11, 13, 'sp4_h_r_23')
// (12, 13, 'sp4_h_r_34')
// (13, 9, 'sp4_h_r_1')
// (13, 13, 'sp4_h_r_47')
// (13, 14, 'neigh_op_tnr_6')
// (13, 14, 'sp4_r_v_b_41')
// (13, 15, 'neigh_op_rgt_6')
// (13, 15, 'sp4_r_v_b_28')
// (13, 15, 'sp4_r_v_b_44')
// (13, 16, 'neigh_op_bnr_6')
// (13, 16, 'sp4_r_v_b_17')
// (13, 16, 'sp4_r_v_b_33')
// (13, 17, 'sp4_r_v_b_20')
// (13, 17, 'sp4_r_v_b_4')
// (13, 18, 'sp4_r_v_b_9')
// (14, 9, 'sp12_h_r_0')
// (14, 9, 'sp12_v_t_23')
// (14, 9, 'sp4_h_r_12')
// (14, 10, 'sp12_v_b_23')
// (14, 11, 'sp12_v_b_20')
// (14, 12, 'sp12_v_b_19')
// (14, 13, 'sp12_v_b_16')
// (14, 13, 'sp4_h_l_47')
// (14, 13, 'sp4_h_r_10')
// (14, 13, 'sp4_h_r_6')
// (14, 13, 'sp4_v_t_41')
// (14, 14, 'local_g0_2')
// (14, 14, 'lutff_global/cen')
// (14, 14, 'neigh_op_top_6')
// (14, 14, 'sp12_v_b_15')
// (14, 14, 'sp4_h_r_2')
// (14, 14, 'sp4_v_b_41')
// (14, 14, 'sp4_v_t_44')
// (14, 15, 'lutff_6/out')
// (14, 15, 'sp12_v_b_12')
// (14, 15, 'sp4_v_b_28')
// (14, 15, 'sp4_v_b_44')
// (14, 16, 'neigh_op_bot_6')
// (14, 16, 'sp12_v_b_11')
// (14, 16, 'sp4_v_b_17')
// (14, 16, 'sp4_v_b_33')
// (14, 17, 'sp12_v_b_8')
// (14, 17, 'sp4_v_b_20')
// (14, 17, 'sp4_v_b_4')
// (14, 18, 'sp12_v_b_7')
// (14, 18, 'sp4_v_b_9')
// (14, 19, 'sp12_v_b_4')
// (14, 20, 'sp12_v_b_3')
// (14, 21, 'sp12_v_b_0')
// (15, 9, 'sp12_h_r_3')
// (15, 9, 'sp4_h_r_25')
// (15, 13, 'local_g1_3')
// (15, 13, 'lutff_global/cen')
// (15, 13, 'sp4_h_r_19')
// (15, 13, 'sp4_h_r_23')
// (15, 14, 'neigh_op_tnl_6')
// (15, 14, 'sp4_h_r_15')
// (15, 15, 'neigh_op_lft_6')
// (15, 16, 'neigh_op_bnl_6')
// (16, 9, 'sp12_h_r_4')
// (16, 9, 'sp4_h_r_36')
// (16, 10, 'sp4_r_v_b_43')
// (16, 11, 'sp4_r_v_b_30')
// (16, 12, 'local_g3_3')
// (16, 12, 'lutff_global/cen')
// (16, 12, 'sp4_r_v_b_19')
// (16, 13, 'local_g2_2')
// (16, 13, 'lutff_global/cen')
// (16, 13, 'sp4_h_r_30')
// (16, 13, 'sp4_h_r_34')
// (16, 13, 'sp4_r_v_b_6')
// (16, 14, 'local_g2_2')
// (16, 14, 'lutff_global/cen')
// (16, 14, 'sp4_h_r_26')
// (17, 9, 'sp12_h_r_7')
// (17, 9, 'sp4_h_l_36')
// (17, 9, 'sp4_v_t_43')
// (17, 10, 'sp4_v_b_43')
// (17, 11, 'sp4_v_b_30')
// (17, 12, 'sp4_v_b_19')
// (17, 13, 'sp4_h_r_43')
// (17, 13, 'sp4_h_r_47')
// (17, 13, 'sp4_v_b_6')
// (17, 14, 'sp4_h_r_39')
// (18, 9, 'sp12_h_r_8')
// (18, 13, 'sp4_h_l_43')
// (18, 13, 'sp4_h_l_47')
// (18, 14, 'sp4_h_l_39')
// (19, 9, 'sp12_h_r_11')
// (20, 9, 'sp12_h_r_12')
// (21, 9, 'sp12_h_r_15')
// (22, 9, 'sp12_h_r_16')
// (23, 9, 'sp12_h_r_19')
// (24, 9, 'sp12_h_r_20')
// (25, 9, 'sp12_h_r_23')
// (26, 9, 'sp12_h_l_23')

reg n322 = 0;
// (10, 13, 'sp4_r_v_b_37')
// (10, 14, 'local_g0_0')
// (10, 14, 'lutff_3/in_1')
// (10, 14, 'sp4_r_v_b_24')
// (10, 15, 'sp4_r_v_b_13')
// (10, 16, 'sp4_r_v_b_0')
// (11, 12, 'sp4_v_t_37')
// (11, 13, 'sp4_v_b_37')
// (11, 14, 'sp4_v_b_24')
// (11, 15, 'sp4_v_b_13')
// (11, 16, 'sp4_h_r_7')
// (11, 16, 'sp4_v_b_0')
// (12, 16, 'sp4_h_r_18')
// (13, 15, 'neigh_op_tnr_5')
// (13, 16, 'neigh_op_rgt_5')
// (13, 16, 'sp4_h_r_31')
// (13, 17, 'neigh_op_bnr_5')
// (14, 15, 'neigh_op_top_5')
// (14, 16, 'local_g1_5')
// (14, 16, 'lutff_5/in_3')
// (14, 16, 'lutff_5/out')
// (14, 16, 'sp4_h_r_42')
// (14, 17, 'neigh_op_bot_5')
// (15, 15, 'neigh_op_tnl_5')
// (15, 16, 'neigh_op_lft_5')
// (15, 16, 'sp4_h_l_42')
// (15, 17, 'neigh_op_bnl_5')

wire n323;
// (10, 14, 'neigh_op_tnr_0')
// (10, 15, 'neigh_op_rgt_0')
// (10, 16, 'neigh_op_bnr_0')
// (11, 14, 'neigh_op_top_0')
// (11, 15, 'lutff_0/out')
// (11, 16, 'neigh_op_bot_0')
// (12, 14, 'neigh_op_tnl_0')
// (12, 15, 'local_g0_0')
// (12, 15, 'lutff_0/in_2')
// (12, 15, 'neigh_op_lft_0')
// (12, 16, 'neigh_op_bnl_0')

wire n324;
// (10, 14, 'neigh_op_tnr_1')
// (10, 15, 'neigh_op_rgt_1')
// (10, 16, 'neigh_op_bnr_1')
// (11, 14, 'neigh_op_top_1')
// (11, 15, 'lutff_1/out')
// (11, 16, 'neigh_op_bot_1')
// (12, 14, 'neigh_op_tnl_1')
// (12, 15, 'local_g0_1')
// (12, 15, 'lutff_1/in_2')
// (12, 15, 'neigh_op_lft_1')
// (12, 16, 'neigh_op_bnl_1')

wire n325;
// (10, 14, 'neigh_op_tnr_2')
// (10, 15, 'neigh_op_rgt_2')
// (10, 16, 'neigh_op_bnr_2')
// (11, 14, 'neigh_op_top_2')
// (11, 15, 'lutff_2/out')
// (11, 16, 'neigh_op_bot_2')
// (12, 14, 'neigh_op_tnl_2')
// (12, 15, 'local_g0_2')
// (12, 15, 'lutff_2/in_2')
// (12, 15, 'neigh_op_lft_2')
// (12, 16, 'neigh_op_bnl_2')

wire n326;
// (10, 14, 'neigh_op_tnr_3')
// (10, 15, 'neigh_op_rgt_3')
// (10, 16, 'neigh_op_bnr_3')
// (11, 14, 'neigh_op_top_3')
// (11, 15, 'lutff_3/out')
// (11, 16, 'neigh_op_bot_3')
// (12, 14, 'neigh_op_tnl_3')
// (12, 15, 'local_g0_3')
// (12, 15, 'lutff_3/in_2')
// (12, 15, 'neigh_op_lft_3')
// (12, 16, 'neigh_op_bnl_3')

wire n327;
// (10, 14, 'neigh_op_tnr_4')
// (10, 15, 'neigh_op_rgt_4')
// (10, 16, 'neigh_op_bnr_4')
// (11, 14, 'neigh_op_top_4')
// (11, 15, 'lutff_4/out')
// (11, 16, 'neigh_op_bot_4')
// (12, 14, 'neigh_op_tnl_4')
// (12, 15, 'local_g0_4')
// (12, 15, 'lutff_4/in_2')
// (12, 15, 'neigh_op_lft_4')
// (12, 16, 'neigh_op_bnl_4')

wire n328;
// (10, 14, 'neigh_op_tnr_5')
// (10, 15, 'neigh_op_rgt_5')
// (10, 16, 'neigh_op_bnr_5')
// (11, 14, 'neigh_op_top_5')
// (11, 15, 'lutff_5/out')
// (11, 16, 'neigh_op_bot_5')
// (12, 14, 'neigh_op_tnl_5')
// (12, 15, 'local_g0_5')
// (12, 15, 'lutff_5/in_2')
// (12, 15, 'neigh_op_lft_5')
// (12, 16, 'neigh_op_bnl_5')

wire n329;
// (10, 14, 'neigh_op_tnr_6')
// (10, 15, 'neigh_op_rgt_6')
// (10, 16, 'neigh_op_bnr_6')
// (11, 14, 'neigh_op_top_6')
// (11, 15, 'lutff_6/out')
// (11, 16, 'neigh_op_bot_6')
// (12, 14, 'neigh_op_tnl_6')
// (12, 15, 'local_g0_6')
// (12, 15, 'lutff_6/in_2')
// (12, 15, 'neigh_op_lft_6')
// (12, 16, 'neigh_op_bnl_6')

wire n330;
// (10, 14, 'neigh_op_tnr_7')
// (10, 15, 'neigh_op_rgt_7')
// (10, 16, 'neigh_op_bnr_7')
// (11, 14, 'neigh_op_top_7')
// (11, 15, 'lutff_7/out')
// (11, 16, 'neigh_op_bot_7')
// (12, 14, 'neigh_op_tnl_7')
// (12, 15, 'local_g0_7')
// (12, 15, 'lutff_7/in_2')
// (12, 15, 'neigh_op_lft_7')
// (12, 16, 'neigh_op_bnl_7')

wire n331;
// (10, 14, 'sp12_h_r_0')
// (11, 14, 'sp12_h_r_3')
// (12, 14, 'sp12_h_r_4')
// (13, 14, 'sp12_h_r_7')
// (14, 14, 'sp12_h_r_8')
// (15, 14, 'sp12_h_r_11')
// (15, 14, 'sp4_h_r_7')
// (16, 14, 'sp12_h_r_12')
// (16, 14, 'sp4_h_r_18')
// (17, 14, 'sp12_h_r_15')
// (17, 14, 'sp4_h_r_31')
// (18, 14, 'sp12_h_r_16')
// (18, 14, 'sp4_h_r_42')
// (18, 15, 'sp4_r_v_b_42')
// (18, 16, 'sp4_r_v_b_31')
// (18, 17, 'sp4_r_v_b_18')
// (18, 18, 'sp4_r_v_b_7')
// (18, 19, 'sp4_r_v_b_47')
// (18, 20, 'sp4_r_v_b_34')
// (18, 21, 'sp4_r_v_b_23')
// (18, 22, 'sp4_r_v_b_10')
// (19, 14, 'sp12_h_r_19')
// (19, 14, 'sp4_h_l_42')
// (19, 14, 'sp4_v_t_42')
// (19, 15, 'sp4_v_b_42')
// (19, 16, 'sp4_v_b_31')
// (19, 17, 'sp4_v_b_18')
// (19, 18, 'sp4_v_b_7')
// (19, 18, 'sp4_v_t_47')
// (19, 19, 'sp4_v_b_47')
// (19, 20, 'sp4_v_b_34')
// (19, 21, 'local_g1_7')
// (19, 21, 'lutff_2/in_0')
// (19, 21, 'sp4_v_b_23')
// (19, 22, 'sp4_v_b_10')
// (20, 14, 'sp12_h_r_20')
// (21, 14, 'sp12_h_r_23')
// (22, 2, 'sp12_h_r_0')
// (22, 2, 'sp12_v_t_23')
// (22, 3, 'sp12_v_b_23')
// (22, 4, 'sp12_v_b_20')
// (22, 5, 'sp12_v_b_19')
// (22, 6, 'sp12_v_b_16')
// (22, 7, 'sp12_v_b_15')
// (22, 8, 'sp12_v_b_12')
// (22, 9, 'sp12_v_b_11')
// (22, 10, 'sp12_v_b_8')
// (22, 11, 'sp12_v_b_7')
// (22, 12, 'sp12_v_b_4')
// (22, 13, 'sp12_v_b_3')
// (22, 14, 'sp12_h_l_23')
// (22, 14, 'sp12_v_b_0')
// (23, 2, 'sp12_h_r_3')
// (24, 2, 'sp12_h_r_4')
// (25, 2, 'sp12_h_r_7')
// (26, 2, 'sp12_h_r_8')
// (27, 2, 'sp12_h_r_11')
// (28, 2, 'sp12_h_r_12')
// (29, 2, 'sp12_h_r_15')
// (30, 2, 'sp12_h_r_16')
// (31, 2, 'sp12_h_r_19')
// (32, 1, 'neigh_op_tnr_2')
// (32, 1, 'neigh_op_tnr_6')
// (32, 2, 'neigh_op_rgt_2')
// (32, 2, 'neigh_op_rgt_6')
// (32, 2, 'sp12_h_r_20')
// (32, 3, 'neigh_op_bnr_2')
// (32, 3, 'neigh_op_bnr_6')
// (33, 2, 'io_1/D_IN_0')
// (33, 2, 'span12_horz_20')

wire n332;
// (10, 15, 'lutff_0/cout')
// (10, 15, 'lutff_1/in_3')

wire n333;
// (10, 15, 'lutff_1/cout')
// (10, 15, 'lutff_2/in_3')

wire n334;
// (10, 15, 'lutff_2/cout')
// (10, 15, 'lutff_3/in_3')

wire n335;
// (10, 15, 'lutff_3/cout')
// (10, 15, 'lutff_4/in_3')

wire n336;
// (10, 15, 'lutff_4/cout')
// (10, 15, 'lutff_5/in_3')

wire n337;
// (10, 15, 'lutff_5/cout')
// (10, 15, 'lutff_6/in_3')

wire n338;
// (10, 15, 'lutff_6/cout')
// (10, 15, 'lutff_7/in_3')

wire n339;
// (10, 15, 'lutff_7/cout')
// (10, 16, 'carry_in')
// (10, 16, 'carry_in_mux')
// (10, 16, 'lutff_0/in_3')

reg n340 = 0;
// (10, 15, 'neigh_op_tnr_3')
// (10, 16, 'neigh_op_rgt_3')
// (10, 17, 'neigh_op_bnr_3')
// (11, 15, 'neigh_op_top_3')
// (11, 16, 'local_g1_3')
// (11, 16, 'lutff_0/in_0')
// (11, 16, 'lutff_3/out')
// (11, 17, 'neigh_op_bot_3')
// (12, 15, 'neigh_op_tnl_3')
// (12, 16, 'local_g0_3')
// (12, 16, 'lutff_5/in_0')
// (12, 16, 'neigh_op_lft_3')
// (12, 17, 'neigh_op_bnl_3')

wire n341;
// (10, 15, 'neigh_op_tnr_4')
// (10, 16, 'neigh_op_rgt_4')
// (10, 17, 'neigh_op_bnr_4')
// (11, 15, 'neigh_op_top_4')
// (11, 16, 'lutff_4/out')
// (11, 17, 'neigh_op_bot_4')
// (12, 15, 'neigh_op_tnl_4')
// (12, 16, 'local_g0_4')
// (12, 16, 'lutff_5/in_1')
// (12, 16, 'neigh_op_lft_4')
// (12, 17, 'neigh_op_bnl_4')

wire n342;
// (10, 15, 'neigh_op_tnr_5')
// (10, 16, 'neigh_op_rgt_5')
// (10, 16, 'sp4_r_v_b_42')
// (10, 17, 'neigh_op_bnr_5')
// (10, 17, 'sp4_r_v_b_31')
// (10, 18, 'sp4_r_v_b_18')
// (10, 19, 'sp4_r_v_b_7')
// (11, 15, 'neigh_op_top_5')
// (11, 15, 'sp4_v_t_42')
// (11, 16, 'local_g1_5')
// (11, 16, 'lutff_1/in_1')
// (11, 16, 'lutff_5/out')
// (11, 16, 'sp4_v_b_42')
// (11, 17, 'local_g3_7')
// (11, 17, 'lutff_1/in_3')
// (11, 17, 'neigh_op_bot_5')
// (11, 17, 'sp4_v_b_31')
// (11, 18, 'sp4_v_b_18')
// (11, 19, 'sp4_v_b_7')
// (12, 15, 'neigh_op_tnl_5')
// (12, 16, 'neigh_op_lft_5')
// (12, 17, 'neigh_op_bnl_5')

reg n343 = 0;
// (10, 15, 'neigh_op_tnr_6')
// (10, 16, 'neigh_op_rgt_6')
// (10, 17, 'neigh_op_bnr_6')
// (11, 15, 'neigh_op_top_6')
// (11, 16, 'local_g3_6')
// (11, 16, 'lutff_4/in_1')
// (11, 16, 'lutff_5/in_2')
// (11, 16, 'lutff_6/out')
// (11, 16, 'lutff_7/in_2')
// (11, 17, 'neigh_op_bot_6')
// (12, 15, 'neigh_op_tnl_6')
// (12, 16, 'neigh_op_lft_6')
// (12, 17, 'neigh_op_bnl_6')

wire n344;
// (10, 15, 'neigh_op_tnr_7')
// (10, 16, 'neigh_op_rgt_7')
// (10, 17, 'neigh_op_bnr_7')
// (11, 15, 'neigh_op_top_7')
// (11, 16, 'lutff_7/out')
// (11, 17, 'local_g0_7')
// (11, 17, 'lutff_5/in_0')
// (11, 17, 'neigh_op_bot_7')
// (12, 15, 'neigh_op_tnl_7')
// (12, 16, 'neigh_op_lft_7')
// (12, 17, 'neigh_op_bnl_7')

reg n345 = 0;
// (10, 15, 'sp4_r_v_b_42')
// (10, 16, 'sp4_r_v_b_31')
// (10, 17, 'sp4_r_v_b_18')
// (10, 18, 'sp4_r_v_b_7')
// (10, 21, 'sp4_h_r_7')
// (11, 14, 'sp4_v_t_42')
// (11, 15, 'sp4_v_b_42')
// (11, 16, 'sp4_v_b_31')
// (11, 17, 'local_g1_2')
// (11, 17, 'lutff_3/in_0')
// (11, 17, 'sp4_v_b_18')
// (11, 18, 'local_g0_7')
// (11, 18, 'lutff_5/in_2')
// (11, 18, 'sp4_h_r_7')
// (11, 18, 'sp4_v_b_7')
// (11, 21, 'sp4_h_r_18')
// (12, 18, 'sp4_h_r_18')
// (12, 21, 'local_g2_7')
// (12, 21, 'lutff_5/in_2')
// (12, 21, 'sp4_h_r_31')
// (13, 17, 'local_g2_5')
// (13, 17, 'local_g3_5')
// (13, 17, 'lutff_0/in_3')
// (13, 17, 'lutff_1/in_1')
// (13, 17, 'neigh_op_tnr_5')
// (13, 18, 'local_g3_5')
// (13, 18, 'lutff_5/in_3')
// (13, 18, 'neigh_op_rgt_5')
// (13, 18, 'sp4_h_r_31')
// (13, 18, 'sp4_r_v_b_42')
// (13, 19, 'neigh_op_bnr_5')
// (13, 19, 'sp4_r_v_b_31')
// (13, 20, 'sp4_r_v_b_18')
// (13, 21, 'sp4_h_r_42')
// (13, 21, 'sp4_r_v_b_7')
// (13, 22, 'local_g2_5')
// (13, 22, 'lutff_5/in_2')
// (13, 22, 'sp4_r_v_b_37')
// (13, 23, 'sp4_r_v_b_24')
// (13, 24, 'sp4_r_v_b_13')
// (13, 25, 'sp4_r_v_b_0')
// (14, 17, 'neigh_op_top_5')
// (14, 17, 'sp4_v_t_42')
// (14, 18, 'local_g1_5')
// (14, 18, 'lutff_5/in_1')
// (14, 18, 'lutff_5/out')
// (14, 18, 'sp4_h_r_42')
// (14, 18, 'sp4_v_b_42')
// (14, 19, 'neigh_op_bot_5')
// (14, 19, 'sp4_r_v_b_42')
// (14, 19, 'sp4_v_b_31')
// (14, 20, 'sp4_r_v_b_31')
// (14, 20, 'sp4_v_b_18')
// (14, 21, 'sp4_h_l_42')
// (14, 21, 'sp4_r_v_b_18')
// (14, 21, 'sp4_v_b_7')
// (14, 21, 'sp4_v_t_37')
// (14, 22, 'sp4_r_v_b_7')
// (14, 22, 'sp4_v_b_37')
// (14, 23, 'sp4_v_b_24')
// (14, 24, 'sp4_v_b_13')
// (14, 25, 'sp4_v_b_0')
// (15, 17, 'neigh_op_tnl_5')
// (15, 18, 'neigh_op_lft_5')
// (15, 18, 'sp4_h_l_42')
// (15, 18, 'sp4_v_t_42')
// (15, 19, 'neigh_op_bnl_5')
// (15, 19, 'sp4_v_b_42')
// (15, 20, 'local_g2_7')
// (15, 20, 'lutff_5/in_2')
// (15, 20, 'sp4_v_b_31')
// (15, 21, 'sp4_v_b_18')
// (15, 22, 'sp4_h_r_1')
// (15, 22, 'sp4_v_b_7')
// (16, 22, 'sp4_h_r_12')
// (17, 22, 'local_g3_1')
// (17, 22, 'lutff_5/in_1')
// (17, 22, 'sp4_h_r_25')
// (18, 22, 'sp4_h_r_36')
// (19, 22, 'sp4_h_l_36')

wire n346;
// (10, 16, 'lutff_0/cout')
// (10, 16, 'lutff_1/in_3')

wire n347;
// (10, 16, 'lutff_1/cout')
// (10, 16, 'lutff_2/in_3')

wire n348;
// (10, 16, 'lutff_2/cout')
// (10, 16, 'lutff_3/in_3')

wire n349;
// (10, 16, 'lutff_3/cout')
// (10, 16, 'lutff_4/in_3')

wire n350;
// (10, 16, 'lutff_4/cout')
// (10, 16, 'lutff_5/in_3')

wire n351;
// (10, 16, 'lutff_5/cout')
// (10, 16, 'lutff_6/in_3')

wire n352;
// (10, 16, 'lutff_6/cout')
// (10, 16, 'lutff_7/in_3')

wire n353;
// (10, 16, 'lutff_7/cout')
// (10, 17, 'carry_in')
// (10, 17, 'carry_in_mux')
// (10, 17, 'lutff_0/in_3')

wire n354;
// (10, 16, 'neigh_op_tnr_3')
// (10, 17, 'neigh_op_rgt_3')
// (10, 17, 'sp4_h_r_11')
// (10, 18, 'neigh_op_bnr_3')
// (11, 16, 'neigh_op_top_3')
// (11, 17, 'lutff_3/out')
// (11, 17, 'sp4_h_r_22')
// (11, 18, 'neigh_op_bot_3')
// (12, 16, 'neigh_op_tnl_3')
// (12, 17, 'neigh_op_lft_3')
// (12, 17, 'sp4_h_r_35')
// (12, 18, 'neigh_op_bnl_3')
// (13, 17, 'sp4_h_r_46')
// (13, 18, 'sp4_r_v_b_41')
// (13, 19, 'sp4_r_v_b_28')
// (13, 20, 'sp4_r_v_b_17')
// (13, 21, 'sp4_r_v_b_4')
// (13, 22, 'sp4_r_v_b_41')
// (13, 23, 'sp4_r_v_b_28')
// (13, 24, 'sp4_r_v_b_17')
// (13, 25, 'local_g1_4')
// (13, 25, 'lutff_0/in_1')
// (13, 25, 'sp4_r_v_b_4')
// (14, 17, 'sp4_h_l_46')
// (14, 17, 'sp4_v_t_41')
// (14, 18, 'sp4_v_b_41')
// (14, 19, 'sp4_v_b_28')
// (14, 20, 'sp4_v_b_17')
// (14, 21, 'sp4_v_b_4')
// (14, 21, 'sp4_v_t_41')
// (14, 22, 'sp4_v_b_41')
// (14, 23, 'sp4_v_b_28')
// (14, 24, 'sp4_v_b_17')
// (14, 25, 'sp4_h_r_4')
// (14, 25, 'sp4_v_b_4')
// (15, 25, 'sp4_h_r_17')
// (16, 25, 'sp4_h_r_28')
// (17, 25, 'local_g2_1')
// (17, 25, 'lutff_0/in_1')
// (17, 25, 'sp4_h_r_41')
// (18, 25, 'sp4_h_l_41')

wire n355;
// (10, 16, 'neigh_op_tnr_4')
// (10, 17, 'neigh_op_rgt_4')
// (10, 18, 'neigh_op_bnr_4')
// (11, 16, 'local_g1_4')
// (11, 16, 'lutff_0/in_1')
// (11, 16, 'lutff_3/in_0')
// (11, 16, 'neigh_op_top_4')
// (11, 17, 'lutff_4/out')
// (11, 18, 'neigh_op_bot_4')
// (12, 16, 'neigh_op_tnl_4')
// (12, 17, 'neigh_op_lft_4')
// (12, 18, 'neigh_op_bnl_4')

wire n356;
// (10, 16, 'neigh_op_tnr_5')
// (10, 17, 'neigh_op_rgt_5')
// (10, 18, 'neigh_op_bnr_5')
// (11, 16, 'neigh_op_top_5')
// (11, 17, 'lutff_5/out')
// (11, 18, 'neigh_op_bot_5')
// (12, 16, 'neigh_op_tnl_5')
// (12, 17, 'local_g0_5')
// (12, 17, 'local_g1_5')
// (12, 17, 'lutff_0/in_2')
// (12, 17, 'lutff_0/in_3')
// (12, 17, 'neigh_op_lft_5')
// (12, 18, 'neigh_op_bnl_5')

wire n357;
// (10, 16, 'neigh_op_tnr_7')
// (10, 17, 'neigh_op_rgt_7')
// (10, 18, 'neigh_op_bnr_7')
// (11, 16, 'local_g1_7')
// (11, 16, 'lutff_1/in_3')
// (11, 16, 'neigh_op_top_7')
// (11, 17, 'lutff_7/out')
// (11, 18, 'neigh_op_bot_7')
// (12, 16, 'neigh_op_tnl_7')
// (12, 17, 'neigh_op_lft_7')
// (12, 18, 'neigh_op_bnl_7')

reg n358 = 0;
// (10, 16, 'sp4_h_r_0')
// (11, 16, 'local_g0_5')
// (11, 16, 'lutff_4/in_3')
// (11, 16, 'lutff_5/in_0')
// (11, 16, 'lutff_6/in_3')
// (11, 16, 'lutff_7/in_0')
// (11, 16, 'sp4_h_r_13')
// (12, 16, 'sp4_h_r_24')
// (13, 13, 'sp4_r_v_b_42')
// (13, 14, 'sp4_r_v_b_31')
// (13, 15, 'sp4_r_v_b_18')
// (13, 16, 'sp4_h_r_37')
// (13, 16, 'sp4_r_v_b_7')
// (14, 11, 'neigh_op_tnr_1')
// (14, 12, 'neigh_op_rgt_1')
// (14, 12, 'sp4_h_r_7')
// (14, 12, 'sp4_v_t_42')
// (14, 13, 'neigh_op_bnr_1')
// (14, 13, 'sp4_v_b_42')
// (14, 14, 'sp4_v_b_31')
// (14, 15, 'local_g0_2')
// (14, 15, 'lutff_7/in_3')
// (14, 15, 'sp4_v_b_18')
// (14, 16, 'sp4_h_l_37')
// (14, 16, 'sp4_v_b_7')
// (15, 11, 'neigh_op_top_1')
// (15, 12, 'local_g3_1')
// (15, 12, 'lutff_1/in_3')
// (15, 12, 'lutff_1/out')
// (15, 12, 'sp4_h_r_18')
// (15, 13, 'neigh_op_bot_1')
// (16, 11, 'neigh_op_tnl_1')
// (16, 12, 'neigh_op_lft_1')
// (16, 12, 'sp4_h_r_31')
// (16, 13, 'neigh_op_bnl_1')
// (17, 12, 'sp4_h_r_42')
// (18, 12, 'sp4_h_l_42')

wire n359;
// (10, 16, 'sp4_r_v_b_38')
// (10, 17, 'sp4_r_v_b_27')
// (10, 18, 'sp4_r_v_b_14')
// (10, 19, 'local_g1_3')
// (10, 19, 'lutff_global/cen')
// (10, 19, 'sp4_r_v_b_3')
// (11, 15, 'sp4_h_r_9')
// (11, 15, 'sp4_v_t_38')
// (11, 16, 'sp4_v_b_38')
// (11, 17, 'sp4_v_b_27')
// (11, 18, 'sp4_v_b_14')
// (11, 19, 'sp4_v_b_3')
// (12, 15, 'sp4_h_r_20')
// (13, 15, 'sp4_h_r_33')
// (14, 12, 'sp4_r_v_b_44')
// (14, 13, 'neigh_op_tnr_2')
// (14, 13, 'sp4_r_v_b_33')
// (14, 14, 'neigh_op_rgt_2')
// (14, 14, 'sp4_r_v_b_20')
// (14, 15, 'neigh_op_bnr_2')
// (14, 15, 'sp4_h_r_44')
// (14, 15, 'sp4_r_v_b_9')
// (15, 11, 'sp4_v_t_44')
// (15, 12, 'sp4_v_b_44')
// (15, 13, 'neigh_op_top_2')
// (15, 13, 'sp4_v_b_33')
// (15, 14, 'lutff_2/out')
// (15, 14, 'sp4_v_b_20')
// (15, 15, 'neigh_op_bot_2')
// (15, 15, 'sp4_h_l_44')
// (15, 15, 'sp4_v_b_9')
// (16, 13, 'neigh_op_tnl_2')
// (16, 14, 'neigh_op_lft_2')
// (16, 15, 'neigh_op_bnl_2')

wire n360;
// (10, 17, 'lutff_0/cout')
// (10, 17, 'lutff_1/in_3')

wire n361;
// (10, 17, 'lutff_1/cout')
// (10, 17, 'lutff_2/in_3')

wire n362;
// (10, 17, 'lutff_2/cout')
// (10, 17, 'lutff_3/in_3')

wire n363;
// (10, 17, 'lutff_3/cout')
// (10, 17, 'lutff_4/in_3')

wire n364;
// (10, 17, 'lutff_4/cout')
// (10, 17, 'lutff_5/in_3')

wire n365;
// (10, 17, 'lutff_7/cout')
// (10, 18, 'carry_in')
// (10, 18, 'carry_in_mux')
// (10, 18, 'lutff_0/in_3')

wire n366;
// (10, 17, 'neigh_op_tnr_0')
// (10, 18, 'neigh_op_rgt_0')
// (10, 19, 'neigh_op_bnr_0')
// (11, 17, 'neigh_op_top_0')
// (11, 18, 'local_g3_0')
// (11, 18, 'lutff_0/in_1')
// (11, 18, 'lutff_0/out')
// (11, 19, 'neigh_op_bot_0')
// (12, 17, 'neigh_op_tnl_0')
// (12, 18, 'neigh_op_lft_0')
// (12, 19, 'neigh_op_bnl_0')

wire n367;
// (10, 17, 'neigh_op_tnr_1')
// (10, 18, 'neigh_op_rgt_1')
// (10, 19, 'neigh_op_bnr_1')
// (11, 17, 'neigh_op_top_1')
// (11, 18, 'local_g1_1')
// (11, 18, 'lutff_1/in_1')
// (11, 18, 'lutff_1/out')
// (11, 19, 'neigh_op_bot_1')
// (12, 17, 'neigh_op_tnl_1')
// (12, 18, 'neigh_op_lft_1')
// (12, 19, 'neigh_op_bnl_1')

wire n368;
// (10, 17, 'neigh_op_tnr_2')
// (10, 18, 'neigh_op_rgt_2')
// (10, 19, 'neigh_op_bnr_2')
// (11, 17, 'neigh_op_top_2')
// (11, 18, 'local_g1_2')
// (11, 18, 'lutff_2/in_1')
// (11, 18, 'lutff_2/out')
// (11, 19, 'neigh_op_bot_2')
// (12, 17, 'neigh_op_tnl_2')
// (12, 18, 'neigh_op_lft_2')
// (12, 19, 'neigh_op_bnl_2')

wire n369;
// (10, 17, 'neigh_op_tnr_3')
// (10, 18, 'neigh_op_rgt_3')
// (10, 19, 'neigh_op_bnr_3')
// (11, 17, 'neigh_op_top_3')
// (11, 18, 'local_g1_3')
// (11, 18, 'lutff_3/in_1')
// (11, 18, 'lutff_3/out')
// (11, 19, 'neigh_op_bot_3')
// (12, 17, 'neigh_op_tnl_3')
// (12, 18, 'neigh_op_lft_3')
// (12, 19, 'neigh_op_bnl_3')

wire n370;
// (10, 17, 'neigh_op_tnr_4')
// (10, 18, 'neigh_op_rgt_4')
// (10, 19, 'neigh_op_bnr_4')
// (11, 17, 'neigh_op_top_4')
// (11, 18, 'local_g1_4')
// (11, 18, 'lutff_4/in_1')
// (11, 18, 'lutff_4/out')
// (11, 19, 'neigh_op_bot_4')
// (12, 17, 'neigh_op_tnl_4')
// (12, 18, 'neigh_op_lft_4')
// (12, 19, 'neigh_op_bnl_4')

wire n371;
// (10, 17, 'neigh_op_tnr_5')
// (10, 18, 'neigh_op_rgt_5')
// (10, 19, 'neigh_op_bnr_5')
// (11, 17, 'neigh_op_top_5')
// (11, 18, 'local_g1_5')
// (11, 18, 'lutff_5/in_1')
// (11, 18, 'lutff_5/out')
// (11, 19, 'neigh_op_bot_5')
// (12, 17, 'neigh_op_tnl_5')
// (12, 18, 'neigh_op_lft_5')
// (12, 19, 'neigh_op_bnl_5')

wire n372;
// (10, 17, 'neigh_op_tnr_6')
// (10, 18, 'neigh_op_rgt_6')
// (10, 19, 'neigh_op_bnr_6')
// (11, 17, 'neigh_op_top_6')
// (11, 18, 'local_g1_6')
// (11, 18, 'lutff_6/in_1')
// (11, 18, 'lutff_6/out')
// (11, 19, 'neigh_op_bot_6')
// (12, 17, 'neigh_op_tnl_6')
// (12, 18, 'neigh_op_lft_6')
// (12, 19, 'neigh_op_bnl_6')

wire n373;
// (10, 17, 'neigh_op_tnr_7')
// (10, 18, 'neigh_op_rgt_7')
// (10, 19, 'neigh_op_bnr_7')
// (11, 17, 'neigh_op_top_7')
// (11, 18, 'local_g1_7')
// (11, 18, 'lutff_7/in_1')
// (11, 18, 'lutff_7/out')
// (11, 19, 'neigh_op_bot_7')
// (12, 17, 'neigh_op_tnl_7')
// (12, 18, 'neigh_op_lft_7')
// (12, 19, 'neigh_op_bnl_7')

wire n374;
// (10, 17, 'sp4_h_r_3')
// (11, 17, 'local_g1_6')
// (11, 17, 'lutff_4/in_1')
// (11, 17, 'lutff_7/in_0')
// (11, 17, 'sp4_h_r_14')
// (12, 16, 'neigh_op_tnr_3')
// (12, 17, 'neigh_op_rgt_3')
// (12, 17, 'sp4_h_r_27')
// (12, 18, 'neigh_op_bnr_3')
// (13, 16, 'neigh_op_top_3')
// (13, 16, 'sp12_v_t_22')
// (13, 17, 'lutff_3/out')
// (13, 17, 'sp12_v_b_22')
// (13, 17, 'sp4_h_r_38')
// (13, 17, 'sp4_h_r_6')
// (13, 18, 'neigh_op_bot_3')
// (13, 18, 'sp12_v_b_21')
// (13, 19, 'sp12_v_b_18')
// (13, 20, 'sp12_v_b_17')
// (13, 21, 'local_g2_6')
// (13, 21, 'lutff_3/in_1')
// (13, 21, 'sp12_v_b_14')
// (13, 22, 'sp12_v_b_13')
// (13, 23, 'sp12_v_b_10')
// (13, 24, 'sp12_v_b_9')
// (13, 25, 'local_g2_6')
// (13, 25, 'lutff_0/in_0')
// (13, 25, 'sp12_v_b_6')
// (13, 26, 'sp12_v_b_5')
// (13, 27, 'sp12_v_b_2')
// (13, 28, 'sp12_v_b_1')
// (14, 16, 'neigh_op_tnl_3')
// (14, 17, 'neigh_op_lft_3')
// (14, 17, 'sp4_h_l_38')
// (14, 17, 'sp4_h_r_19')
// (14, 18, 'neigh_op_bnl_3')
// (15, 17, 'sp4_h_r_30')
// (16, 17, 'sp4_h_r_43')
// (16, 18, 'sp4_r_v_b_46')
// (16, 19, 'sp4_r_v_b_35')
// (16, 20, 'sp4_r_v_b_22')
// (16, 21, 'sp4_r_v_b_11')
// (16, 22, 'sp4_r_v_b_46')
// (16, 23, 'sp4_r_v_b_35')
// (16, 24, 'sp4_r_v_b_22')
// (16, 25, 'sp4_r_v_b_11')
// (17, 17, 'sp4_h_l_43')
// (17, 17, 'sp4_v_t_46')
// (17, 18, 'sp4_v_b_46')
// (17, 19, 'sp4_v_b_35')
// (17, 20, 'sp4_v_b_22')
// (17, 21, 'sp4_v_b_11')
// (17, 21, 'sp4_v_t_46')
// (17, 22, 'sp4_v_b_46')
// (17, 23, 'sp4_v_b_35')
// (17, 24, 'sp4_v_b_22')
// (17, 25, 'local_g1_3')
// (17, 25, 'lutff_0/in_2')
// (17, 25, 'sp4_v_b_11')

wire n375;
// (10, 18, 'neigh_op_tnr_0')
// (10, 19, 'neigh_op_rgt_0')
// (10, 20, 'neigh_op_bnr_0')
// (11, 18, 'neigh_op_top_0')
// (11, 19, 'local_g3_0')
// (11, 19, 'lutff_0/in_1')
// (11, 19, 'lutff_0/out')
// (11, 20, 'neigh_op_bot_0')
// (12, 18, 'neigh_op_tnl_0')
// (12, 19, 'neigh_op_lft_0')
// (12, 20, 'neigh_op_bnl_0')

wire n376;
// (10, 18, 'neigh_op_tnr_1')
// (10, 19, 'neigh_op_rgt_1')
// (10, 20, 'neigh_op_bnr_1')
// (11, 18, 'neigh_op_top_1')
// (11, 19, 'local_g3_1')
// (11, 19, 'lutff_1/in_1')
// (11, 19, 'lutff_1/out')
// (11, 20, 'neigh_op_bot_1')
// (12, 18, 'neigh_op_tnl_1')
// (12, 19, 'neigh_op_lft_1')
// (12, 20, 'neigh_op_bnl_1')

wire n377;
// (10, 18, 'neigh_op_tnr_2')
// (10, 19, 'neigh_op_rgt_2')
// (10, 20, 'neigh_op_bnr_2')
// (11, 18, 'neigh_op_top_2')
// (11, 19, 'local_g1_2')
// (11, 19, 'lutff_2/in_1')
// (11, 19, 'lutff_2/out')
// (11, 20, 'neigh_op_bot_2')
// (12, 18, 'neigh_op_tnl_2')
// (12, 19, 'neigh_op_lft_2')
// (12, 20, 'neigh_op_bnl_2')

wire n378;
// (10, 18, 'neigh_op_tnr_3')
// (10, 19, 'neigh_op_rgt_3')
// (10, 20, 'neigh_op_bnr_3')
// (11, 18, 'neigh_op_top_3')
// (11, 19, 'local_g1_3')
// (11, 19, 'lutff_3/in_1')
// (11, 19, 'lutff_3/out')
// (11, 20, 'neigh_op_bot_3')
// (12, 18, 'neigh_op_tnl_3')
// (12, 19, 'neigh_op_lft_3')
// (12, 20, 'neigh_op_bnl_3')

wire n379;
// (10, 18, 'neigh_op_tnr_4')
// (10, 19, 'neigh_op_rgt_4')
// (10, 20, 'neigh_op_bnr_4')
// (11, 18, 'neigh_op_top_4')
// (11, 19, 'local_g3_4')
// (11, 19, 'lutff_4/in_1')
// (11, 19, 'lutff_4/out')
// (11, 20, 'neigh_op_bot_4')
// (12, 18, 'neigh_op_tnl_4')
// (12, 19, 'neigh_op_lft_4')
// (12, 20, 'neigh_op_bnl_4')

wire n380;
// (10, 18, 'neigh_op_tnr_5')
// (10, 19, 'neigh_op_rgt_5')
// (10, 20, 'neigh_op_bnr_5')
// (11, 18, 'neigh_op_top_5')
// (11, 19, 'local_g1_5')
// (11, 19, 'lutff_5/in_1')
// (11, 19, 'lutff_5/out')
// (11, 20, 'neigh_op_bot_5')
// (12, 18, 'neigh_op_tnl_5')
// (12, 19, 'neigh_op_lft_5')
// (12, 20, 'neigh_op_bnl_5')

wire n381;
// (10, 18, 'neigh_op_tnr_6')
// (10, 19, 'neigh_op_rgt_6')
// (10, 20, 'neigh_op_bnr_6')
// (11, 18, 'neigh_op_top_6')
// (11, 19, 'local_g1_6')
// (11, 19, 'lutff_6/in_1')
// (11, 19, 'lutff_6/out')
// (11, 20, 'neigh_op_bot_6')
// (12, 18, 'neigh_op_tnl_6')
// (12, 19, 'neigh_op_lft_6')
// (12, 20, 'neigh_op_bnl_6')

wire n382;
// (10, 18, 'neigh_op_tnr_7')
// (10, 19, 'neigh_op_rgt_7')
// (10, 20, 'neigh_op_bnr_7')
// (11, 18, 'neigh_op_top_7')
// (11, 19, 'local_g1_7')
// (11, 19, 'lutff_7/in_1')
// (11, 19, 'lutff_7/out')
// (11, 20, 'neigh_op_bot_7')
// (12, 18, 'neigh_op_tnl_7')
// (12, 19, 'neigh_op_lft_7')
// (12, 20, 'neigh_op_bnl_7')

wire n383;
// (10, 18, 'sp12_h_r_0')
// (11, 18, 'sp12_h_r_3')
// (12, 18, 'sp12_h_r_4')
// (13, 18, 'sp12_h_r_7')
// (14, 18, 'sp12_h_r_8')
// (15, 18, 'sp12_h_r_11')
// (16, 18, 'sp12_h_r_12')
// (17, 18, 'sp12_h_r_15')
// (18, 18, 'sp12_h_r_16')
// (18, 19, 'sp4_r_v_b_46')
// (18, 20, 'sp4_r_v_b_35')
// (18, 21, 'sp4_r_v_b_22')
// (18, 22, 'sp4_r_v_b_11')
// (19, 18, 'sp12_h_r_19')
// (19, 18, 'sp4_h_r_11')
// (19, 18, 'sp4_v_t_46')
// (19, 19, 'sp4_v_b_46')
// (19, 20, 'sp4_v_b_35')
// (19, 21, 'local_g0_6')
// (19, 21, 'lutff_0/in_2')
// (19, 21, 'sp4_v_b_22')
// (19, 22, 'sp4_v_b_11')
// (20, 18, 'sp12_h_r_20')
// (20, 18, 'sp4_h_r_22')
// (21, 18, 'sp12_h_r_23')
// (21, 18, 'sp4_h_r_35')
// (22, 6, 'sp12_h_r_0')
// (22, 6, 'sp12_v_t_23')
// (22, 7, 'sp12_v_b_23')
// (22, 8, 'sp12_v_b_20')
// (22, 9, 'sp12_v_b_19')
// (22, 10, 'sp12_v_b_16')
// (22, 11, 'sp12_v_b_15')
// (22, 12, 'sp12_v_b_12')
// (22, 13, 'sp12_v_b_11')
// (22, 14, 'sp12_v_b_8')
// (22, 15, 'sp12_v_b_7')
// (22, 16, 'sp12_v_b_4')
// (22, 17, 'sp12_v_b_3')
// (22, 18, 'sp12_h_l_23')
// (22, 18, 'sp12_v_b_0')
// (22, 18, 'sp4_h_r_46')
// (23, 6, 'sp12_h_r_3')
// (23, 18, 'sp4_h_l_46')
// (24, 6, 'sp12_h_r_4')
// (25, 6, 'sp12_h_r_7')
// (26, 6, 'sp12_h_r_8')
// (27, 6, 'sp12_h_r_11')
// (28, 6, 'sp12_h_r_12')
// (29, 6, 'sp12_h_r_15')
// (30, 6, 'sp12_h_r_16')
// (31, 6, 'sp12_h_r_19')
// (32, 5, 'neigh_op_tnr_2')
// (32, 5, 'neigh_op_tnr_6')
// (32, 6, 'neigh_op_rgt_2')
// (32, 6, 'neigh_op_rgt_6')
// (32, 6, 'sp12_h_r_20')
// (32, 7, 'neigh_op_bnr_2')
// (32, 7, 'neigh_op_bnr_6')
// (33, 6, 'io_1/D_IN_0')
// (33, 6, 'span12_horz_20')

wire n384;
// (10, 18, 'sp12_h_r_1')
// (11, 18, 'sp12_h_r_2')
// (12, 17, 'neigh_op_tnr_7')
// (12, 18, 'neigh_op_rgt_7')
// (12, 18, 'sp12_h_r_5')
// (12, 19, 'neigh_op_bnr_7')
// (13, 17, 'neigh_op_top_7')
// (13, 18, 'local_g0_7')
// (13, 18, 'lutff_7/in_2')
// (13, 18, 'lutff_7/out')
// (13, 18, 'sp12_h_r_6')
// (13, 19, 'neigh_op_bot_7')
// (14, 17, 'neigh_op_tnl_7')
// (14, 18, 'neigh_op_lft_7')
// (14, 18, 'sp12_h_r_9')
// (14, 19, 'neigh_op_bnl_7')
// (15, 18, 'sp12_h_r_10')
// (16, 18, 'sp12_h_r_13')
// (17, 18, 'local_g1_6')
// (17, 18, 'lutff_7/in_2')
// (17, 18, 'sp12_h_r_14')
// (18, 18, 'sp12_h_r_17')
// (19, 18, 'sp12_h_r_18')
// (20, 18, 'sp12_h_r_21')
// (21, 18, 'sp12_h_r_22')
// (22, 18, 'sp12_h_l_22')

reg n385 = 0;
// (10, 18, 'sp4_h_r_3')
// (11, 15, 'sp4_r_v_b_36')
// (11, 16, 'sp4_r_v_b_25')
// (11, 17, 'local_g2_4')
// (11, 17, 'lutff_6/in_0')
// (11, 17, 'sp4_r_v_b_12')
// (11, 18, 'local_g0_6')
// (11, 18, 'lutff_0/in_2')
// (11, 18, 'sp4_h_r_14')
// (11, 18, 'sp4_r_v_b_1')
// (11, 19, 'sp4_r_v_b_36')
// (11, 20, 'sp4_r_v_b_25')
// (11, 21, 'sp4_r_v_b_12')
// (11, 22, 'sp4_r_v_b_1')
// (12, 14, 'sp4_v_t_36')
// (12, 15, 'sp4_v_b_36')
// (12, 16, 'sp4_v_b_25')
// (12, 17, 'sp4_v_b_12')
// (12, 18, 'sp4_h_r_27')
// (12, 18, 'sp4_h_r_8')
// (12, 18, 'sp4_v_b_1')
// (12, 18, 'sp4_v_t_36')
// (12, 19, 'sp4_v_b_36')
// (12, 20, 'sp4_v_b_25')
// (12, 21, 'local_g0_4')
// (12, 21, 'lutff_0/in_2')
// (12, 21, 'sp4_v_b_12')
// (12, 22, 'sp4_v_b_1')
// (13, 17, 'local_g2_0')
// (13, 17, 'lutff_5/in_3')
// (13, 17, 'lutff_7/in_3')
// (13, 17, 'neigh_op_tnr_0')
// (13, 18, 'local_g3_0')
// (13, 18, 'lutff_0/in_3')
// (13, 18, 'neigh_op_rgt_0')
// (13, 18, 'sp4_h_r_21')
// (13, 18, 'sp4_h_r_38')
// (13, 19, 'neigh_op_bnr_0')
// (13, 19, 'sp4_r_v_b_37')
// (13, 20, 'sp4_r_v_b_24')
// (13, 21, 'sp4_r_v_b_13')
// (13, 22, 'local_g1_0')
// (13, 22, 'lutff_0/in_1')
// (13, 22, 'sp4_r_v_b_0')
// (14, 17, 'neigh_op_top_0')
// (14, 17, 'sp4_r_v_b_44')
// (14, 18, 'local_g3_0')
// (14, 18, 'lutff_0/in_1')
// (14, 18, 'lutff_0/out')
// (14, 18, 'sp4_h_l_38')
// (14, 18, 'sp4_h_r_0')
// (14, 18, 'sp4_h_r_32')
// (14, 18, 'sp4_r_v_b_33')
// (14, 18, 'sp4_v_t_37')
// (14, 19, 'neigh_op_bot_0')
// (14, 19, 'sp4_r_v_b_20')
// (14, 19, 'sp4_v_b_37')
// (14, 20, 'sp4_r_v_b_9')
// (14, 20, 'sp4_v_b_24')
// (14, 21, 'sp4_v_b_13')
// (14, 22, 'sp4_v_b_0')
// (15, 16, 'sp4_v_t_44')
// (15, 17, 'neigh_op_tnl_0')
// (15, 17, 'sp4_v_b_44')
// (15, 18, 'neigh_op_lft_0')
// (15, 18, 'sp4_h_r_13')
// (15, 18, 'sp4_h_r_45')
// (15, 18, 'sp4_v_b_33')
// (15, 19, 'neigh_op_bnl_0')
// (15, 19, 'sp4_v_b_20')
// (15, 20, 'local_g1_1')
// (15, 20, 'lutff_0/in_2')
// (15, 20, 'sp4_v_b_9')
// (16, 18, 'sp4_h_l_45')
// (16, 18, 'sp4_h_r_24')
// (17, 18, 'sp4_h_r_37')
// (17, 19, 'sp4_r_v_b_40')
// (17, 20, 'sp4_r_v_b_29')
// (17, 21, 'sp4_r_v_b_16')
// (17, 22, 'local_g1_5')
// (17, 22, 'lutff_0/in_2')
// (17, 22, 'sp4_r_v_b_5')
// (18, 18, 'sp4_h_l_37')
// (18, 18, 'sp4_v_t_40')
// (18, 19, 'sp4_v_b_40')
// (18, 20, 'sp4_v_b_29')
// (18, 21, 'sp4_v_b_16')
// (18, 22, 'sp4_v_b_5')

reg n386 = 0;
// (10, 18, 'sp4_h_r_7')
// (11, 18, 'local_g0_2')
// (11, 18, 'lutff_2/in_2')
// (11, 18, 'sp4_h_r_18')
// (11, 21, 'sp4_h_r_5')
// (12, 18, 'sp4_h_r_31')
// (12, 21, 'local_g1_0')
// (12, 21, 'lutff_2/in_1')
// (12, 21, 'sp4_h_r_16')
// (13, 17, 'local_g3_2')
// (13, 17, 'lutff_6/in_1')
// (13, 17, 'lutff_7/in_2')
// (13, 17, 'neigh_op_tnr_2')
// (13, 18, 'local_g3_2')
// (13, 18, 'lutff_2/in_3')
// (13, 18, 'neigh_op_rgt_2')
// (13, 18, 'sp4_h_r_42')
// (13, 19, 'neigh_op_bnr_2')
// (13, 19, 'sp4_r_v_b_42')
// (13, 20, 'sp4_r_v_b_31')
// (13, 21, 'sp4_h_r_29')
// (13, 21, 'sp4_r_v_b_18')
// (13, 22, 'local_g1_7')
// (13, 22, 'lutff_2/in_2')
// (13, 22, 'sp4_r_v_b_7')
// (14, 17, 'neigh_op_top_2')
// (14, 18, 'local_g1_2')
// (14, 18, 'lutff_2/in_1')
// (14, 18, 'lutff_2/out')
// (14, 18, 'sp4_h_l_42')
// (14, 18, 'sp4_h_r_4')
// (14, 18, 'sp4_r_v_b_37')
// (14, 18, 'sp4_v_t_42')
// (14, 19, 'neigh_op_bot_2')
// (14, 19, 'sp4_r_v_b_24')
// (14, 19, 'sp4_v_b_42')
// (14, 20, 'sp4_r_v_b_13')
// (14, 20, 'sp4_v_b_31')
// (14, 21, 'sp4_h_r_40')
// (14, 21, 'sp4_r_v_b_0')
// (14, 21, 'sp4_v_b_18')
// (14, 22, 'sp4_v_b_7')
// (15, 17, 'neigh_op_tnl_2')
// (15, 17, 'sp4_v_t_37')
// (15, 18, 'neigh_op_lft_2')
// (15, 18, 'sp4_h_r_17')
// (15, 18, 'sp4_v_b_37')
// (15, 19, 'neigh_op_bnl_2')
// (15, 19, 'sp4_v_b_24')
// (15, 20, 'local_g1_5')
// (15, 20, 'lutff_2/in_2')
// (15, 20, 'sp4_v_b_13')
// (15, 21, 'sp4_h_l_40')
// (15, 21, 'sp4_v_b_0')
// (16, 18, 'sp4_h_r_28')
// (17, 18, 'sp4_h_r_41')
// (17, 19, 'sp4_r_v_b_44')
// (17, 20, 'sp4_r_v_b_33')
// (17, 21, 'sp4_r_v_b_20')
// (17, 22, 'local_g2_1')
// (17, 22, 'lutff_2/in_1')
// (17, 22, 'sp4_r_v_b_9')
// (18, 18, 'sp4_h_l_41')
// (18, 18, 'sp4_v_t_44')
// (18, 19, 'sp4_v_b_44')
// (18, 20, 'sp4_v_b_33')
// (18, 21, 'sp4_v_b_20')
// (18, 22, 'sp4_v_b_9')

wire n387;
// (10, 19, 'neigh_op_tnr_0')
// (10, 20, 'neigh_op_rgt_0')
// (10, 21, 'neigh_op_bnr_0')
// (11, 19, 'neigh_op_top_0')
// (11, 20, 'local_g3_0')
// (11, 20, 'lutff_0/in_1')
// (11, 20, 'lutff_0/out')
// (11, 21, 'neigh_op_bot_0')
// (12, 19, 'neigh_op_tnl_0')
// (12, 20, 'neigh_op_lft_0')
// (12, 21, 'neigh_op_bnl_0')

wire n388;
// (10, 19, 'neigh_op_tnr_1')
// (10, 20, 'neigh_op_rgt_1')
// (10, 21, 'neigh_op_bnr_1')
// (11, 19, 'neigh_op_top_1')
// (11, 20, 'local_g3_1')
// (11, 20, 'lutff_1/in_1')
// (11, 20, 'lutff_1/out')
// (11, 21, 'neigh_op_bot_1')
// (12, 19, 'neigh_op_tnl_1')
// (12, 20, 'neigh_op_lft_1')
// (12, 21, 'neigh_op_bnl_1')

wire n389;
// (10, 19, 'neigh_op_tnr_2')
// (10, 20, 'neigh_op_rgt_2')
// (10, 21, 'neigh_op_bnr_2')
// (11, 19, 'neigh_op_top_2')
// (11, 20, 'local_g1_2')
// (11, 20, 'lutff_2/in_1')
// (11, 20, 'lutff_2/out')
// (11, 21, 'neigh_op_bot_2')
// (12, 19, 'neigh_op_tnl_2')
// (12, 20, 'neigh_op_lft_2')
// (12, 21, 'neigh_op_bnl_2')

wire n390;
// (10, 19, 'neigh_op_tnr_3')
// (10, 20, 'neigh_op_rgt_3')
// (10, 21, 'neigh_op_bnr_3')
// (11, 19, 'neigh_op_top_3')
// (11, 20, 'local_g1_3')
// (11, 20, 'lutff_3/in_1')
// (11, 20, 'lutff_3/out')
// (11, 21, 'neigh_op_bot_3')
// (12, 19, 'neigh_op_tnl_3')
// (12, 20, 'neigh_op_lft_3')
// (12, 21, 'neigh_op_bnl_3')

wire n391;
// (10, 19, 'neigh_op_tnr_4')
// (10, 20, 'neigh_op_rgt_4')
// (10, 21, 'neigh_op_bnr_4')
// (11, 19, 'neigh_op_top_4')
// (11, 20, 'local_g3_4')
// (11, 20, 'lutff_4/in_1')
// (11, 20, 'lutff_4/out')
// (11, 21, 'neigh_op_bot_4')
// (12, 19, 'neigh_op_tnl_4')
// (12, 20, 'neigh_op_lft_4')
// (12, 21, 'neigh_op_bnl_4')

wire n392;
// (10, 19, 'neigh_op_tnr_5')
// (10, 20, 'neigh_op_rgt_5')
// (10, 21, 'neigh_op_bnr_5')
// (11, 19, 'neigh_op_top_5')
// (11, 20, 'local_g1_5')
// (11, 20, 'lutff_5/in_1')
// (11, 20, 'lutff_5/out')
// (11, 21, 'neigh_op_bot_5')
// (12, 19, 'neigh_op_tnl_5')
// (12, 20, 'neigh_op_lft_5')
// (12, 21, 'neigh_op_bnl_5')

wire n393;
// (10, 19, 'neigh_op_tnr_6')
// (10, 20, 'neigh_op_rgt_6')
// (10, 21, 'neigh_op_bnr_6')
// (11, 19, 'neigh_op_top_6')
// (11, 20, 'local_g1_6')
// (11, 20, 'lutff_6/in_1')
// (11, 20, 'lutff_6/out')
// (11, 21, 'neigh_op_bot_6')
// (12, 19, 'neigh_op_tnl_6')
// (12, 20, 'neigh_op_lft_6')
// (12, 21, 'neigh_op_bnl_6')

wire n394;
// (10, 19, 'neigh_op_tnr_7')
// (10, 20, 'neigh_op_rgt_7')
// (10, 21, 'neigh_op_bnr_7')
// (11, 19, 'neigh_op_top_7')
// (11, 20, 'local_g1_7')
// (11, 20, 'lutff_7/in_1')
// (11, 20, 'lutff_7/out')
// (11, 21, 'neigh_op_bot_7')
// (12, 19, 'neigh_op_tnl_7')
// (12, 20, 'neigh_op_lft_7')
// (12, 21, 'neigh_op_bnl_7')

wire n395;
// (10, 19, 'sp12_h_r_1')
// (11, 19, 'sp12_h_r_2')
// (12, 18, 'neigh_op_tnr_7')
// (12, 19, 'neigh_op_rgt_7')
// (12, 19, 'sp12_h_r_5')
// (12, 20, 'neigh_op_bnr_7')
// (13, 18, 'neigh_op_top_7')
// (13, 19, 'local_g1_7')
// (13, 19, 'lutff_7/in_1')
// (13, 19, 'lutff_7/out')
// (13, 19, 'sp12_h_r_6')
// (13, 20, 'neigh_op_bot_7')
// (14, 18, 'neigh_op_tnl_7')
// (14, 19, 'neigh_op_lft_7')
// (14, 19, 'sp12_h_r_9')
// (14, 20, 'neigh_op_bnl_7')
// (15, 19, 'sp12_h_r_10')
// (16, 19, 'sp12_h_r_13')
// (17, 19, 'local_g1_6')
// (17, 19, 'lutff_7/in_2')
// (17, 19, 'sp12_h_r_14')
// (18, 19, 'sp12_h_r_17')
// (19, 19, 'sp12_h_r_18')
// (20, 19, 'sp12_h_r_21')
// (21, 19, 'sp12_h_r_22')
// (22, 19, 'sp12_h_l_22')

reg n396 = 0;
// (10, 20, 'sp4_h_r_1')
// (11, 20, 'local_g1_4')
// (11, 20, 'lutff_5/in_2')
// (11, 20, 'sp4_h_r_12')
// (11, 23, 'sp4_h_r_6')
// (12, 20, 'sp4_h_r_25')
// (12, 23, 'local_g1_3')
// (12, 23, 'lutff_5/in_1')
// (12, 23, 'sp4_h_r_19')
// (13, 17, 'sp4_r_v_b_47')
// (13, 18, 'sp4_r_v_b_34')
// (13, 19, 'neigh_op_tnr_5')
// (13, 19, 'sp4_r_v_b_23')
// (13, 20, 'local_g3_5')
// (13, 20, 'lutff_5/in_3')
// (13, 20, 'neigh_op_rgt_5')
// (13, 20, 'sp4_h_r_36')
// (13, 20, 'sp4_r_v_b_10')
// (13, 21, 'neigh_op_bnr_5')
// (13, 21, 'sp4_r_v_b_47')
// (13, 22, 'sp4_r_v_b_34')
// (13, 23, 'sp4_h_r_30')
// (13, 23, 'sp4_r_v_b_23')
// (13, 24, 'local_g2_2')
// (13, 24, 'lutff_5/in_1')
// (13, 24, 'sp4_r_v_b_10')
// (14, 16, 'sp4_v_t_47')
// (14, 17, 'local_g2_7')
// (14, 17, 'lutff_1/in_0')
// (14, 17, 'sp4_v_b_47')
// (14, 18, 'sp4_v_b_34')
// (14, 19, 'neigh_op_top_5')
// (14, 19, 'sp4_v_b_23')
// (14, 20, 'local_g1_5')
// (14, 20, 'lutff_5/in_1')
// (14, 20, 'lutff_5/out')
// (14, 20, 'sp4_h_l_36')
// (14, 20, 'sp4_h_r_10')
// (14, 20, 'sp4_r_v_b_43')
// (14, 20, 'sp4_v_b_10')
// (14, 20, 'sp4_v_t_47')
// (14, 21, 'neigh_op_bot_5')
// (14, 21, 'sp4_r_v_b_30')
// (14, 21, 'sp4_v_b_47')
// (14, 22, 'sp4_r_v_b_19')
// (14, 22, 'sp4_v_b_34')
// (14, 23, 'sp4_h_r_43')
// (14, 23, 'sp4_r_v_b_6')
// (14, 23, 'sp4_v_b_23')
// (14, 24, 'sp4_v_b_10')
// (15, 19, 'neigh_op_tnl_5')
// (15, 19, 'sp4_v_t_43')
// (15, 20, 'neigh_op_lft_5')
// (15, 20, 'sp4_h_r_23')
// (15, 20, 'sp4_v_b_43')
// (15, 21, 'neigh_op_bnl_5')
// (15, 21, 'sp4_v_b_30')
// (15, 22, 'local_g0_3')
// (15, 22, 'lutff_5/in_2')
// (15, 22, 'sp4_v_b_19')
// (15, 23, 'sp4_h_l_43')
// (15, 23, 'sp4_v_b_6')
// (16, 20, 'sp4_h_r_34')
// (17, 20, 'local_g2_7')
// (17, 20, 'lutff_5/in_0')
// (17, 20, 'sp4_h_r_47')
// (17, 21, 'sp4_r_v_b_38')
// (17, 22, 'sp4_r_v_b_27')
// (17, 23, 'sp4_r_v_b_14')
// (17, 24, 'local_g1_3')
// (17, 24, 'lutff_5/in_1')
// (17, 24, 'sp4_r_v_b_3')
// (18, 20, 'sp4_h_l_47')
// (18, 20, 'sp4_v_t_38')
// (18, 21, 'sp4_v_b_38')
// (18, 22, 'sp4_v_b_27')
// (18, 23, 'sp4_v_b_14')
// (18, 24, 'sp4_v_b_3')

reg n397 = 0;
// (10, 20, 'sp4_h_r_2')
// (11, 20, 'local_g0_7')
// (11, 20, 'lutff_1/in_2')
// (11, 20, 'sp4_h_r_15')
// (11, 21, 'sp4_r_v_b_41')
// (11, 22, 'sp4_r_v_b_28')
// (11, 23, 'sp4_r_v_b_17')
// (11, 24, 'sp4_r_v_b_4')
// (12, 20, 'sp4_h_r_10')
// (12, 20, 'sp4_h_r_26')
// (12, 20, 'sp4_v_t_41')
// (12, 21, 'sp4_v_b_41')
// (12, 22, 'sp4_v_b_28')
// (12, 23, 'local_g1_1')
// (12, 23, 'lutff_1/in_1')
// (12, 23, 'sp4_v_b_17')
// (12, 24, 'sp4_h_r_4')
// (12, 24, 'sp4_v_b_4')
// (13, 17, 'sp4_r_v_b_39')
// (13, 18, 'sp4_r_v_b_26')
// (13, 19, 'neigh_op_tnr_1')
// (13, 19, 'sp4_r_v_b_15')
// (13, 20, 'local_g2_1')
// (13, 20, 'lutff_1/in_0')
// (13, 20, 'neigh_op_rgt_1')
// (13, 20, 'sp4_h_r_23')
// (13, 20, 'sp4_h_r_39')
// (13, 20, 'sp4_r_v_b_2')
// (13, 21, 'neigh_op_bnr_1')
// (13, 24, 'local_g1_1')
// (13, 24, 'lutff_1/in_1')
// (13, 24, 'sp4_h_r_17')
// (14, 16, 'sp4_v_t_39')
// (14, 17, 'local_g3_7')
// (14, 17, 'lutff_1/in_3')
// (14, 17, 'sp4_v_b_39')
// (14, 18, 'sp4_v_b_26')
// (14, 19, 'neigh_op_top_1')
// (14, 19, 'sp4_r_v_b_46')
// (14, 19, 'sp4_v_b_15')
// (14, 20, 'local_g3_1')
// (14, 20, 'lutff_1/in_1')
// (14, 20, 'lutff_1/out')
// (14, 20, 'sp4_h_l_39')
// (14, 20, 'sp4_h_r_2')
// (14, 20, 'sp4_h_r_34')
// (14, 20, 'sp4_r_v_b_35')
// (14, 20, 'sp4_v_b_2')
// (14, 21, 'neigh_op_bot_1')
// (14, 21, 'sp4_r_v_b_22')
// (14, 22, 'sp4_r_v_b_11')
// (14, 24, 'sp4_h_r_28')
// (15, 18, 'sp4_v_t_46')
// (15, 19, 'neigh_op_tnl_1')
// (15, 19, 'sp4_v_b_46')
// (15, 20, 'neigh_op_lft_1')
// (15, 20, 'sp4_h_r_15')
// (15, 20, 'sp4_h_r_47')
// (15, 20, 'sp4_v_b_35')
// (15, 21, 'neigh_op_bnl_1')
// (15, 21, 'sp4_v_b_22')
// (15, 22, 'local_g1_3')
// (15, 22, 'lutff_1/in_1')
// (15, 22, 'sp4_v_b_11')
// (15, 24, 'sp4_h_r_41')
// (16, 20, 'sp4_h_l_47')
// (16, 20, 'sp4_h_r_26')
// (16, 24, 'sp4_h_l_41')
// (17, 20, 'local_g3_7')
// (17, 20, 'lutff_1/in_3')
// (17, 20, 'sp4_h_r_39')
// (17, 21, 'sp4_r_v_b_42')
// (17, 22, 'sp4_r_v_b_31')
// (17, 23, 'sp4_r_v_b_18')
// (17, 24, 'local_g1_7')
// (17, 24, 'lutff_1/in_1')
// (17, 24, 'sp4_r_v_b_7')
// (18, 20, 'sp4_h_l_39')
// (18, 20, 'sp4_v_t_42')
// (18, 21, 'sp4_v_b_42')
// (18, 22, 'sp4_v_b_31')
// (18, 23, 'sp4_v_b_18')
// (18, 24, 'sp4_v_b_7')

reg n398 = 0;
// (10, 20, 'sp4_h_r_3')
// (11, 20, 'local_g0_6')
// (11, 20, 'lutff_0/in_2')
// (11, 20, 'sp4_h_r_14')
// (11, 21, 'sp4_r_v_b_45')
// (11, 22, 'sp4_r_v_b_32')
// (11, 23, 'sp4_r_v_b_21')
// (11, 24, 'sp4_r_v_b_8')
// (12, 20, 'sp4_h_r_27')
// (12, 20, 'sp4_h_r_8')
// (12, 20, 'sp4_v_t_45')
// (12, 21, 'sp4_v_b_45')
// (12, 22, 'sp4_v_b_32')
// (12, 23, 'local_g1_5')
// (12, 23, 'lutff_0/in_2')
// (12, 23, 'sp4_v_b_21')
// (12, 24, 'sp4_h_r_2')
// (12, 24, 'sp4_v_b_8')
// (13, 17, 'sp4_r_v_b_37')
// (13, 18, 'sp4_r_v_b_24')
// (13, 19, 'neigh_op_tnr_0')
// (13, 19, 'sp4_r_v_b_13')
// (13, 20, 'local_g3_0')
// (13, 20, 'lutff_0/in_3')
// (13, 20, 'neigh_op_rgt_0')
// (13, 20, 'sp4_h_r_21')
// (13, 20, 'sp4_h_r_38')
// (13, 20, 'sp4_r_v_b_0')
// (13, 21, 'neigh_op_bnr_0')
// (13, 24, 'local_g1_7')
// (13, 24, 'lutff_0/in_2')
// (13, 24, 'sp4_h_r_15')
// (14, 16, 'sp4_v_t_37')
// (14, 17, 'local_g2_5')
// (14, 17, 'lutff_0/in_3')
// (14, 17, 'sp4_v_b_37')
// (14, 18, 'sp4_v_b_24')
// (14, 19, 'neigh_op_top_0')
// (14, 19, 'sp4_r_v_b_44')
// (14, 19, 'sp4_v_b_13')
// (14, 20, 'local_g3_0')
// (14, 20, 'lutff_0/in_1')
// (14, 20, 'lutff_0/out')
// (14, 20, 'sp4_h_l_38')
// (14, 20, 'sp4_h_r_0')
// (14, 20, 'sp4_h_r_32')
// (14, 20, 'sp4_r_v_b_33')
// (14, 20, 'sp4_v_b_0')
// (14, 21, 'neigh_op_bot_0')
// (14, 21, 'sp4_r_v_b_20')
// (14, 22, 'sp4_r_v_b_9')
// (14, 24, 'sp4_h_r_26')
// (15, 18, 'sp4_v_t_44')
// (15, 19, 'neigh_op_tnl_0')
// (15, 19, 'sp4_v_b_44')
// (15, 20, 'neigh_op_lft_0')
// (15, 20, 'sp4_h_r_13')
// (15, 20, 'sp4_h_r_45')
// (15, 20, 'sp4_v_b_33')
// (15, 21, 'neigh_op_bnl_0')
// (15, 21, 'sp4_v_b_20')
// (15, 22, 'local_g0_1')
// (15, 22, 'lutff_0/in_1')
// (15, 22, 'sp4_v_b_9')
// (15, 24, 'sp4_h_r_39')
// (16, 20, 'sp4_h_l_45')
// (16, 20, 'sp4_h_r_24')
// (16, 24, 'sp4_h_l_39')
// (17, 20, 'local_g2_5')
// (17, 20, 'lutff_0/in_3')
// (17, 20, 'sp4_h_r_37')
// (17, 21, 'sp4_r_v_b_37')
// (17, 22, 'sp4_r_v_b_24')
// (17, 23, 'sp4_r_v_b_13')
// (17, 24, 'local_g1_0')
// (17, 24, 'lutff_0/in_1')
// (17, 24, 'sp4_r_v_b_0')
// (18, 20, 'sp4_h_l_37')
// (18, 20, 'sp4_v_t_37')
// (18, 21, 'sp4_v_b_37')
// (18, 22, 'sp4_v_b_24')
// (18, 23, 'sp4_v_b_13')
// (18, 24, 'sp4_v_b_0')

reg n399 = 0;
// (10, 21, 'neigh_op_tnr_1')
// (10, 22, 'neigh_op_rgt_1')
// (10, 22, 'sp4_h_r_7')
// (10, 23, 'neigh_op_bnr_1')
// (11, 21, 'neigh_op_top_1')
// (11, 22, 'lutff_1/out')
// (11, 22, 'sp4_h_r_18')
// (11, 23, 'neigh_op_bot_1')
// (12, 21, 'neigh_op_tnl_1')
// (12, 22, 'neigh_op_lft_1')
// (12, 22, 'sp4_h_r_31')
// (12, 23, 'neigh_op_bnl_1')
// (13, 22, 'local_g3_2')
// (13, 22, 'lutff_1/in_0')
// (13, 22, 'sp4_h_r_42')
// (14, 22, 'sp4_h_l_42')

reg n400 = 0;
// (10, 21, 'neigh_op_tnr_2')
// (10, 22, 'neigh_op_rgt_2')
// (10, 22, 'sp4_h_r_9')
// (10, 23, 'neigh_op_bnr_2')
// (11, 21, 'neigh_op_top_2')
// (11, 22, 'lutff_2/out')
// (11, 22, 'sp4_h_r_20')
// (11, 23, 'neigh_op_bot_2')
// (12, 21, 'neigh_op_tnl_2')
// (12, 22, 'neigh_op_lft_2')
// (12, 22, 'sp4_h_r_33')
// (12, 23, 'neigh_op_bnl_2')
// (13, 22, 'local_g3_4')
// (13, 22, 'lutff_2/in_3')
// (13, 22, 'sp4_h_r_44')
// (14, 22, 'sp4_h_l_44')

reg n401 = 0;
// (10, 21, 'neigh_op_tnr_3')
// (10, 22, 'neigh_op_rgt_3')
// (10, 22, 'sp4_h_r_11')
// (10, 23, 'neigh_op_bnr_3')
// (11, 21, 'neigh_op_top_3')
// (11, 22, 'lutff_3/out')
// (11, 22, 'sp4_h_r_22')
// (11, 23, 'neigh_op_bot_3')
// (12, 21, 'neigh_op_tnl_3')
// (12, 22, 'neigh_op_lft_3')
// (12, 22, 'sp4_h_r_35')
// (12, 23, 'neigh_op_bnl_3')
// (13, 22, 'local_g3_6')
// (13, 22, 'lutff_6/in_3')
// (13, 22, 'sp4_h_r_46')
// (14, 22, 'sp4_h_l_46')

reg n402 = 0;
// (10, 21, 'neigh_op_tnr_4')
// (10, 22, 'neigh_op_rgt_4')
// (10, 23, 'neigh_op_bnr_4')
// (11, 21, 'neigh_op_top_4')
// (11, 22, 'lutff_4/out')
// (11, 22, 'sp4_h_r_8')
// (11, 23, 'neigh_op_bot_4')
// (12, 21, 'neigh_op_tnl_4')
// (12, 22, 'neigh_op_lft_4')
// (12, 22, 'sp4_h_r_21')
// (12, 23, 'neigh_op_bnl_4')
// (13, 22, 'local_g3_0')
// (13, 22, 'lutff_4/in_3')
// (13, 22, 'sp4_h_r_32')
// (14, 22, 'sp4_h_r_45')
// (15, 22, 'sp4_h_l_45')

reg n403 = 0;
// (10, 21, 'neigh_op_tnr_5')
// (10, 22, 'neigh_op_rgt_5')
// (10, 22, 'sp12_h_r_1')
// (10, 23, 'neigh_op_bnr_5')
// (11, 21, 'neigh_op_top_5')
// (11, 22, 'lutff_5/out')
// (11, 22, 'sp12_h_r_2')
// (11, 23, 'neigh_op_bot_5')
// (12, 21, 'neigh_op_tnl_5')
// (12, 22, 'neigh_op_lft_5')
// (12, 22, 'sp12_h_r_5')
// (12, 23, 'neigh_op_bnl_5')
// (13, 22, 'local_g0_6')
// (13, 22, 'lutff_5/in_3')
// (13, 22, 'sp12_h_r_6')
// (14, 22, 'sp12_h_r_9')
// (15, 22, 'sp12_h_r_10')
// (16, 22, 'sp12_h_r_13')
// (17, 22, 'sp12_h_r_14')
// (18, 22, 'sp12_h_r_17')
// (19, 22, 'sp12_h_r_18')
// (20, 22, 'sp12_h_r_21')
// (21, 22, 'sp12_h_r_22')
// (22, 22, 'sp12_h_l_22')

reg n404 = 0;
// (10, 21, 'neigh_op_tnr_7')
// (10, 22, 'neigh_op_rgt_7')
// (10, 22, 'sp4_h_r_3')
// (10, 23, 'neigh_op_bnr_7')
// (11, 21, 'neigh_op_top_7')
// (11, 22, 'lutff_7/out')
// (11, 22, 'sp4_h_r_14')
// (11, 23, 'neigh_op_bot_7')
// (12, 21, 'neigh_op_tnl_7')
// (12, 22, 'neigh_op_lft_7')
// (12, 22, 'sp4_h_r_27')
// (12, 23, 'neigh_op_bnl_7')
// (13, 22, 'local_g2_6')
// (13, 22, 'lutff_3/in_3')
// (13, 22, 'sp4_h_r_38')
// (14, 22, 'sp4_h_l_38')

reg io_33_4_1 = 0;
// (10, 21, 'sp12_h_r_0')
// (11, 21, 'sp12_h_r_3')
// (12, 21, 'sp12_h_r_4')
// (13, 21, 'sp12_h_r_7')
// (14, 21, 'sp12_h_r_8')
// (15, 21, 'sp12_h_r_11')
// (16, 21, 'sp12_h_r_12')
// (17, 20, 'neigh_op_tnr_4')
// (17, 21, 'neigh_op_rgt_4')
// (17, 21, 'sp12_h_r_15')
// (17, 22, 'neigh_op_bnr_4')
// (18, 20, 'neigh_op_top_4')
// (18, 21, 'lutff_4/out')
// (18, 21, 'sp12_h_r_16')
// (18, 22, 'neigh_op_bot_4')
// (19, 20, 'neigh_op_tnl_4')
// (19, 21, 'neigh_op_lft_4')
// (19, 21, 'sp12_h_r_19')
// (19, 22, 'neigh_op_bnl_4')
// (20, 21, 'sp12_h_r_20')
// (21, 21, 'sp12_h_r_23')
// (22, 9, 'sp12_h_r_0')
// (22, 9, 'sp12_v_t_23')
// (22, 10, 'sp12_v_b_23')
// (22, 11, 'sp12_v_b_20')
// (22, 12, 'sp12_v_b_19')
// (22, 13, 'sp12_v_b_16')
// (22, 14, 'sp12_v_b_15')
// (22, 15, 'sp12_v_b_12')
// (22, 16, 'sp12_v_b_11')
// (22, 17, 'sp12_v_b_8')
// (22, 18, 'sp12_v_b_7')
// (22, 19, 'sp12_v_b_4')
// (22, 20, 'sp12_v_b_3')
// (22, 21, 'sp12_h_l_23')
// (22, 21, 'sp12_v_b_0')
// (23, 9, 'sp12_h_r_3')
// (24, 9, 'sp12_h_r_4')
// (25, 9, 'sp12_h_r_7')
// (26, 9, 'sp12_h_r_8')
// (27, 9, 'sp12_h_r_11')
// (27, 9, 'sp4_h_r_7')
// (28, 9, 'sp12_h_r_12')
// (28, 9, 'sp4_h_r_18')
// (29, 9, 'sp12_h_r_15')
// (29, 9, 'sp4_h_r_31')
// (30, 6, 'sp4_r_v_b_36')
// (30, 7, 'sp4_r_v_b_25')
// (30, 8, 'sp4_r_v_b_12')
// (30, 9, 'sp12_h_r_16')
// (30, 9, 'sp4_h_r_42')
// (30, 9, 'sp4_r_v_b_1')
// (31, 5, 'sp4_h_r_6')
// (31, 5, 'sp4_v_t_36')
// (31, 6, 'sp4_v_b_36')
// (31, 7, 'sp4_v_b_25')
// (31, 8, 'sp4_v_b_12')
// (31, 9, 'sp12_h_r_19')
// (31, 9, 'sp4_h_l_42')
// (31, 9, 'sp4_v_b_1')
// (32, 5, 'sp4_h_r_19')
// (32, 9, 'sp12_h_r_20')
// (33, 1, 'span4_vert_t_15')
// (33, 2, 'span4_vert_b_15')
// (33, 3, 'span4_vert_b_11')
// (33, 4, 'io_1/D_OUT_0')
// (33, 4, 'io_1/PAD')
// (33, 4, 'local_g0_7')
// (33, 4, 'span4_vert_b_7')
// (33, 5, 'span4_horz_19')
// (33, 5, 'span4_vert_b_3')
// (33, 9, 'span12_horz_20')

wire n406;
// (11, 8, 'neigh_op_tnr_3')
// (11, 9, 'local_g1_3')
// (11, 9, 'lutff_1/in_1')
// (11, 9, 'neigh_op_rgt_3')
// (11, 9, 'sp4_h_r_11')
// (11, 10, 'neigh_op_bnr_3')
// (12, 8, 'neigh_op_top_3')
// (12, 9, 'lutff_3/out')
// (12, 9, 'sp4_h_r_22')
// (12, 10, 'neigh_op_bot_3')
// (13, 8, 'neigh_op_tnl_3')
// (13, 9, 'neigh_op_lft_3')
// (13, 9, 'sp4_h_r_35')
// (13, 10, 'neigh_op_bnl_3')
// (14, 9, 'sp4_h_r_46')
// (15, 9, 'sp4_h_l_46')

wire n407;
// (11, 9, 'lutff_3/lout')
// (11, 9, 'lutff_4/in_2')

wire n408;
// (11, 9, 'lutff_6/lout')
// (11, 9, 'lutff_7/in_2')

wire n409;
// (11, 9, 'neigh_op_tnr_3')
// (11, 10, 'local_g3_3')
// (11, 10, 'lutff_5/in_1')
// (11, 10, 'neigh_op_rgt_3')
// (11, 11, 'neigh_op_bnr_3')
// (12, 9, 'neigh_op_top_3')
// (12, 10, 'lutff_3/out')
// (12, 11, 'neigh_op_bot_3')
// (13, 9, 'neigh_op_tnl_3')
// (13, 10, 'neigh_op_lft_3')
// (13, 11, 'neigh_op_bnl_3')

wire n410;
// (11, 9, 'neigh_op_tnr_7')
// (11, 10, 'neigh_op_rgt_7')
// (11, 11, 'neigh_op_bnr_7')
// (12, 9, 'neigh_op_top_7')
// (12, 10, 'local_g0_7')
// (12, 10, 'lutff_2/in_1')
// (12, 10, 'lutff_7/out')
// (12, 11, 'neigh_op_bot_7')
// (13, 9, 'neigh_op_tnl_7')
// (13, 10, 'neigh_op_lft_7')
// (13, 11, 'neigh_op_bnl_7')

wire n411;
// (11, 10, 'local_g2_7')
// (11, 10, 'lutff_5/in_0')
// (11, 10, 'sp4_r_v_b_39')
// (11, 11, 'sp4_r_v_b_26')
// (11, 12, 'sp4_r_v_b_15')
// (11, 13, 'sp4_r_v_b_2')
// (12, 9, 'sp4_h_r_2')
// (12, 9, 'sp4_v_t_39')
// (12, 10, 'sp4_v_b_39')
// (12, 11, 'sp4_v_b_26')
// (12, 12, 'sp4_v_b_15')
// (12, 13, 'sp4_v_b_2')
// (13, 8, 'neigh_op_tnr_5')
// (13, 9, 'neigh_op_rgt_5')
// (13, 9, 'sp4_h_r_15')
// (13, 10, 'neigh_op_bnr_5')
// (14, 8, 'neigh_op_top_5')
// (14, 9, 'lutff_5/out')
// (14, 9, 'sp4_h_r_26')
// (14, 10, 'neigh_op_bot_5')
// (15, 8, 'neigh_op_tnl_5')
// (15, 9, 'neigh_op_lft_5')
// (15, 9, 'sp4_h_r_39')
// (15, 10, 'neigh_op_bnl_5')
// (16, 9, 'sp4_h_l_39')

wire n412;
// (11, 10, 'lutff_0/lout')
// (11, 10, 'lutff_1/in_2')

wire n413;
// (11, 10, 'lutff_2/lout')
// (11, 10, 'lutff_3/in_2')

reg n414 = 0;
// (11, 10, 'sp12_h_r_0')
// (12, 10, 'sp12_h_r_3')
// (13, 10, 'sp12_h_r_4')
// (14, 10, 'local_g0_7')
// (14, 10, 'lutff_1/in_0')
// (14, 10, 'sp12_h_r_7')
// (15, 10, 'sp12_h_r_8')
// (16, 9, 'neigh_op_tnr_2')
// (16, 10, 'neigh_op_rgt_2')
// (16, 10, 'sp12_h_r_11')
// (16, 11, 'neigh_op_bnr_2')
// (17, 9, 'neigh_op_top_2')
// (17, 10, 'lutff_2/out')
// (17, 10, 'sp12_h_r_12')
// (17, 11, 'neigh_op_bot_2')
// (18, 9, 'neigh_op_tnl_2')
// (18, 10, 'neigh_op_lft_2')
// (18, 10, 'sp12_h_r_15')
// (18, 11, 'neigh_op_bnl_2')
// (19, 10, 'sp12_h_r_16')
// (20, 10, 'sp12_h_r_19')
// (21, 10, 'sp12_h_r_20')
// (22, 10, 'sp12_h_r_23')
// (23, 10, 'sp12_h_l_23')

wire n415;
// (11, 11, 'carry_in_mux')
// (11, 11, 'lutff_0/in_3')

wire n416;
// (11, 11, 'lutff_0/cout')
// (11, 11, 'lutff_1/in_3')

wire n417;
// (11, 11, 'lutff_1/cout')
// (11, 11, 'lutff_2/in_3')

wire n418;
// (11, 11, 'lutff_2/cout')
// (11, 11, 'lutff_3/in_3')

wire n419;
// (11, 11, 'lutff_3/cout')
// (11, 11, 'lutff_4/in_3')

wire n420;
// (11, 11, 'lutff_4/cout')
// (11, 11, 'lutff_5/in_3')

wire n421;
// (11, 11, 'lutff_5/cout')
// (11, 11, 'lutff_6/in_3')

wire n422;
// (11, 11, 'lutff_6/cout')
// (11, 11, 'lutff_7/in_3')

reg n423 = 0;
// (11, 11, 'neigh_op_tnr_0')
// (11, 12, 'local_g3_0')
// (11, 12, 'lutff_6/in_3')
// (11, 12, 'neigh_op_rgt_0')
// (11, 13, 'neigh_op_bnr_0')
// (12, 11, 'neigh_op_top_0')
// (12, 12, 'local_g1_0')
// (12, 12, 'lutff_0/out')
// (12, 12, 'lutff_6/in_3')
// (12, 13, 'neigh_op_bot_0')
// (13, 11, 'neigh_op_tnl_0')
// (13, 12, 'neigh_op_lft_0')
// (13, 13, 'neigh_op_bnl_0')

reg n424 = 0;
// (11, 11, 'neigh_op_tnr_1')
// (11, 12, 'local_g2_1')
// (11, 12, 'lutff_4/in_3')
// (11, 12, 'neigh_op_rgt_1')
// (11, 13, 'neigh_op_bnr_1')
// (12, 11, 'neigh_op_top_1')
// (12, 12, 'local_g3_1')
// (12, 12, 'lutff_1/out')
// (12, 12, 'lutff_7/in_3')
// (12, 13, 'neigh_op_bot_1')
// (13, 11, 'neigh_op_tnl_1')
// (13, 12, 'neigh_op_lft_1')
// (13, 13, 'neigh_op_bnl_1')

reg n425 = 0;
// (11, 11, 'neigh_op_tnr_2')
// (11, 12, 'local_g2_2')
// (11, 12, 'lutff_1/in_3')
// (11, 12, 'neigh_op_rgt_2')
// (11, 13, 'neigh_op_bnr_2')
// (12, 11, 'neigh_op_top_2')
// (12, 12, 'lutff_2/out')
// (12, 13, 'neigh_op_bot_2')
// (13, 11, 'neigh_op_tnl_2')
// (13, 12, 'neigh_op_lft_2')
// (13, 13, 'local_g3_2')
// (13, 13, 'lutff_6/in_3')
// (13, 13, 'neigh_op_bnl_2')

reg n426 = 0;
// (11, 11, 'neigh_op_tnr_3')
// (11, 12, 'local_g3_3')
// (11, 12, 'lutff_0/in_0')
// (11, 12, 'neigh_op_rgt_3')
// (11, 13, 'neigh_op_bnr_3')
// (12, 11, 'neigh_op_top_3')
// (12, 12, 'local_g0_3')
// (12, 12, 'lutff_2/in_3')
// (12, 12, 'lutff_3/out')
// (12, 13, 'neigh_op_bot_3')
// (13, 11, 'neigh_op_tnl_3')
// (13, 12, 'neigh_op_lft_3')
// (13, 13, 'neigh_op_bnl_3')

reg n427 = 0;
// (11, 11, 'neigh_op_tnr_4')
// (11, 12, 'local_g3_4')
// (11, 12, 'lutff_3/in_0')
// (11, 12, 'neigh_op_rgt_4')
// (11, 13, 'neigh_op_bnr_4')
// (12, 11, 'neigh_op_top_4')
// (12, 12, 'local_g0_4')
// (12, 12, 'lutff_1/in_3')
// (12, 12, 'lutff_4/out')
// (12, 13, 'neigh_op_bot_4')
// (13, 11, 'neigh_op_tnl_4')
// (13, 12, 'neigh_op_lft_4')
// (13, 13, 'neigh_op_bnl_4')

reg n428 = 0;
// (11, 11, 'neigh_op_tnr_6')
// (11, 12, 'local_g2_6')
// (11, 12, 'lutff_7/in_3')
// (11, 12, 'neigh_op_rgt_6')
// (11, 13, 'neigh_op_bnr_6')
// (12, 11, 'neigh_op_top_6')
// (12, 12, 'lutff_6/out')
// (12, 13, 'neigh_op_bot_6')
// (13, 11, 'neigh_op_tnl_6')
// (13, 12, 'neigh_op_lft_6')
// (13, 13, 'neigh_op_bnl_6')

reg n429 = 0;
// (11, 11, 'neigh_op_tnr_7')
// (11, 12, 'local_g3_7')
// (11, 12, 'lutff_5/in_3')
// (11, 12, 'neigh_op_rgt_7')
// (11, 13, 'neigh_op_bnr_7')
// (12, 11, 'neigh_op_top_7')
// (12, 12, 'local_g2_7')
// (12, 12, 'lutff_0/in_3')
// (12, 12, 'lutff_7/out')
// (12, 13, 'neigh_op_bot_7')
// (13, 11, 'neigh_op_tnl_7')
// (13, 12, 'neigh_op_lft_7')
// (13, 13, 'neigh_op_bnl_7')

reg n430 = 0;
// (11, 11, 'sp12_h_r_0')
// (12, 11, 'sp12_h_r_3')
// (13, 11, 'sp12_h_r_4')
// (14, 11, 'sp12_h_r_7')
// (15, 11, 'sp12_h_r_8')
// (16, 11, 'sp12_h_r_11')
// (17, 11, 'local_g1_4')
// (17, 11, 'lutff_3/in_0')
// (17, 11, 'sp12_h_r_12')
// (18, 11, 'sp12_h_r_15')
// (19, 11, 'sp12_h_r_16')
// (20, 10, 'neigh_op_tnr_6')
// (20, 11, 'neigh_op_rgt_6')
// (20, 11, 'sp12_h_r_19')
// (20, 12, 'neigh_op_bnr_6')
// (21, 10, 'neigh_op_top_6')
// (21, 11, 'lutff_6/out')
// (21, 11, 'sp12_h_r_20')
// (21, 12, 'neigh_op_bot_6')
// (22, 10, 'neigh_op_tnl_6')
// (22, 11, 'neigh_op_lft_6')
// (22, 11, 'sp12_h_r_23')
// (22, 12, 'neigh_op_bnl_6')
// (23, 11, 'sp12_h_l_23')

reg n431 = 0;
// (11, 12, 'neigh_op_tnr_0')
// (11, 13, 'neigh_op_rgt_0')
// (11, 14, 'local_g0_0')
// (11, 14, 'lutff_0/in_2')
// (11, 14, 'neigh_op_bnr_0')
// (12, 12, 'neigh_op_top_0')
// (12, 13, 'lutff_0/out')
// (12, 14, 'neigh_op_bot_0')
// (13, 12, 'neigh_op_tnl_0')
// (13, 13, 'local_g0_0')
// (13, 13, 'lutff_3/in_1')
// (13, 13, 'neigh_op_lft_0')
// (13, 14, 'neigh_op_bnl_0')

reg n432 = 0;
// (11, 12, 'neigh_op_tnr_1')
// (11, 13, 'neigh_op_rgt_1')
// (11, 14, 'local_g0_1')
// (11, 14, 'lutff_1/in_2')
// (11, 14, 'neigh_op_bnr_1')
// (12, 12, 'neigh_op_top_1')
// (12, 13, 'lutff_1/out')
// (12, 14, 'neigh_op_bot_1')
// (13, 12, 'neigh_op_tnl_1')
// (13, 13, 'neigh_op_lft_1')
// (13, 14, 'neigh_op_bnl_1')

reg n433 = 0;
// (11, 12, 'neigh_op_tnr_2')
// (11, 13, 'neigh_op_rgt_2')
// (11, 14, 'local_g0_2')
// (11, 14, 'lutff_2/in_2')
// (11, 14, 'neigh_op_bnr_2')
// (12, 12, 'neigh_op_top_2')
// (12, 13, 'lutff_2/out')
// (12, 14, 'neigh_op_bot_2')
// (13, 12, 'neigh_op_tnl_2')
// (13, 13, 'neigh_op_lft_2')
// (13, 14, 'neigh_op_bnl_2')

reg n434 = 0;
// (11, 12, 'neigh_op_tnr_3')
// (11, 13, 'neigh_op_rgt_3')
// (11, 14, 'local_g0_3')
// (11, 14, 'lutff_3/in_2')
// (11, 14, 'neigh_op_bnr_3')
// (12, 12, 'neigh_op_top_3')
// (12, 13, 'lutff_3/out')
// (12, 14, 'neigh_op_bot_3')
// (13, 12, 'neigh_op_tnl_3')
// (13, 13, 'neigh_op_lft_3')
// (13, 14, 'neigh_op_bnl_3')

reg n435 = 0;
// (11, 12, 'neigh_op_tnr_4')
// (11, 13, 'neigh_op_rgt_4')
// (11, 14, 'local_g0_4')
// (11, 14, 'lutff_4/in_2')
// (11, 14, 'neigh_op_bnr_4')
// (12, 12, 'neigh_op_top_4')
// (12, 13, 'lutff_4/out')
// (12, 14, 'neigh_op_bot_4')
// (13, 12, 'neigh_op_tnl_4')
// (13, 13, 'neigh_op_lft_4')
// (13, 14, 'neigh_op_bnl_4')

reg n436 = 0;
// (11, 12, 'neigh_op_tnr_5')
// (11, 13, 'neigh_op_rgt_5')
// (11, 14, 'local_g0_5')
// (11, 14, 'lutff_5/in_2')
// (11, 14, 'neigh_op_bnr_5')
// (12, 12, 'neigh_op_top_5')
// (12, 13, 'lutff_5/out')
// (12, 14, 'neigh_op_bot_5')
// (13, 12, 'neigh_op_tnl_5')
// (13, 13, 'neigh_op_lft_5')
// (13, 14, 'neigh_op_bnl_5')

reg n437 = 0;
// (11, 12, 'neigh_op_tnr_6')
// (11, 13, 'neigh_op_rgt_6')
// (11, 14, 'local_g0_6')
// (11, 14, 'lutff_6/in_2')
// (11, 14, 'neigh_op_bnr_6')
// (12, 12, 'neigh_op_top_6')
// (12, 13, 'lutff_6/out')
// (12, 14, 'neigh_op_bot_6')
// (13, 12, 'neigh_op_tnl_6')
// (13, 13, 'neigh_op_lft_6')
// (13, 14, 'neigh_op_bnl_6')

reg n438 = 0;
// (11, 12, 'neigh_op_tnr_7')
// (11, 13, 'neigh_op_rgt_7')
// (11, 14, 'local_g0_7')
// (11, 14, 'lutff_7/in_2')
// (11, 14, 'neigh_op_bnr_7')
// (12, 12, 'neigh_op_top_7')
// (12, 13, 'lutff_7/out')
// (12, 14, 'neigh_op_bot_7')
// (13, 12, 'neigh_op_tnl_7')
// (13, 13, 'neigh_op_lft_7')
// (13, 14, 'neigh_op_bnl_7')

reg n439 = 0;
// (11, 12, 'sp12_h_r_0')
// (12, 12, 'sp12_h_r_3')
// (13, 12, 'sp12_h_r_4')
// (14, 12, 'sp12_h_r_7')
// (15, 12, 'sp12_h_r_8')
// (16, 12, 'sp12_h_r_11')
// (17, 12, 'local_g0_4')
// (17, 12, 'lutff_5/in_3')
// (17, 12, 'sp12_h_r_12')
// (18, 12, 'sp12_h_r_15')
// (19, 12, 'sp12_h_r_16')
// (20, 12, 'sp12_h_r_19')
// (21, 12, 'sp12_h_r_20')
// (22, 12, 'sp12_h_r_23')
// (22, 15, 'neigh_op_tnr_0')
// (22, 16, 'neigh_op_rgt_0')
// (22, 17, 'neigh_op_bnr_0')
// (23, 12, 'sp12_h_l_23')
// (23, 12, 'sp12_v_t_23')
// (23, 13, 'sp12_v_b_23')
// (23, 14, 'sp12_v_b_20')
// (23, 15, 'neigh_op_top_0')
// (23, 15, 'sp12_v_b_19')
// (23, 16, 'lutff_0/out')
// (23, 16, 'sp12_v_b_16')
// (23, 17, 'neigh_op_bot_0')
// (23, 17, 'sp12_v_b_15')
// (23, 18, 'sp12_v_b_12')
// (23, 19, 'sp12_v_b_11')
// (23, 20, 'sp12_v_b_8')
// (23, 21, 'sp12_v_b_7')
// (23, 22, 'sp12_v_b_4')
// (23, 23, 'sp12_v_b_3')
// (23, 24, 'sp12_v_b_0')
// (24, 15, 'neigh_op_tnl_0')
// (24, 16, 'neigh_op_lft_0')
// (24, 17, 'neigh_op_bnl_0')

reg n440 = 0;
// (11, 12, 'sp12_h_r_1')
// (12, 12, 'sp12_h_r_2')
// (13, 12, 'sp12_h_r_5')
// (14, 12, 'sp12_h_r_6')
// (15, 11, 'neigh_op_tnr_1')
// (15, 12, 'neigh_op_rgt_1')
// (15, 12, 'sp12_h_r_9')
// (15, 13, 'neigh_op_bnr_1')
// (15, 15, 'sp4_r_v_b_40')
// (15, 16, 'local_g1_5')
// (15, 16, 'lutff_6/in_0')
// (15, 16, 'sp4_r_v_b_29')
// (15, 17, 'sp4_r_v_b_16')
// (15, 18, 'sp4_r_v_b_5')
// (16, 9, 'sp12_v_t_22')
// (16, 10, 'sp12_v_b_22')
// (16, 11, 'neigh_op_top_1')
// (16, 11, 'sp12_v_b_21')
// (16, 12, 'local_g0_1')
// (16, 12, 'lutff_0/in_1')
// (16, 12, 'lutff_1/out')
// (16, 12, 'lutff_6/in_1')
// (16, 12, 'sp12_h_r_10')
// (16, 12, 'sp12_v_b_18')
// (16, 13, 'local_g0_1')
// (16, 13, 'lutff_2/in_1')
// (16, 13, 'lutff_4/in_1')
// (16, 13, 'lutff_6/in_1')
// (16, 13, 'neigh_op_bot_1')
// (16, 13, 'sp12_v_b_17')
// (16, 14, 'sp12_v_b_14')
// (16, 14, 'sp4_v_t_40')
// (16, 15, 'local_g2_5')
// (16, 15, 'lutff_6/in_3')
// (16, 15, 'sp12_v_b_13')
// (16, 15, 'sp4_v_b_40')
// (16, 16, 'sp12_v_b_10')
// (16, 16, 'sp4_v_b_29')
// (16, 17, 'sp12_v_b_9')
// (16, 17, 'sp4_v_b_16')
// (16, 18, 'sp12_v_b_6')
// (16, 18, 'sp4_v_b_5')
// (16, 19, 'sp12_v_b_5')
// (16, 20, 'sp12_v_b_2')
// (16, 21, 'sp12_v_b_1')
// (17, 11, 'neigh_op_tnl_1')
// (17, 12, 'neigh_op_lft_1')
// (17, 12, 'sp12_h_r_13')
// (17, 13, 'neigh_op_bnl_1')
// (18, 12, 'sp12_h_r_14')
// (19, 12, 'local_g1_1')
// (19, 12, 'lutff_6/in_0')
// (19, 12, 'sp12_h_r_17')
// (20, 12, 'sp12_h_r_18')
// (21, 12, 'sp12_h_r_21')
// (22, 12, 'sp12_h_r_22')
// (23, 12, 'sp12_h_l_22')

wire n441;
// (11, 13, 'local_g0_2')
// (11, 13, 'lutff_global/cen')
// (11, 13, 'sp4_h_r_10')
// (12, 13, 'sp4_h_r_23')
// (13, 13, 'sp4_h_r_34')
// (14, 10, 'sp4_r_v_b_41')
// (14, 11, 'sp4_r_v_b_28')
// (14, 12, 'neigh_op_tnr_2')
// (14, 12, 'sp4_r_v_b_17')
// (14, 13, 'neigh_op_rgt_2')
// (14, 13, 'sp4_h_r_47')
// (14, 13, 'sp4_r_v_b_4')
// (14, 14, 'neigh_op_bnr_2')
// (15, 9, 'sp4_v_t_41')
// (15, 10, 'sp4_v_b_41')
// (15, 11, 'sp4_v_b_28')
// (15, 12, 'neigh_op_top_2')
// (15, 12, 'sp4_v_b_17')
// (15, 13, 'lutff_2/out')
// (15, 13, 'sp4_h_l_47')
// (15, 13, 'sp4_h_r_10')
// (15, 13, 'sp4_v_b_4')
// (15, 14, 'neigh_op_bot_2')
// (16, 12, 'neigh_op_tnl_2')
// (16, 13, 'neigh_op_lft_2')
// (16, 13, 'sp4_h_r_23')
// (16, 14, 'neigh_op_bnl_2')
// (17, 13, 'sp4_h_r_34')
// (18, 13, 'sp4_h_r_47')
// (19, 13, 'sp4_h_l_47')

wire n442;
// (11, 13, 'neigh_op_tnr_0')
// (11, 14, 'neigh_op_rgt_0')
// (11, 15, 'neigh_op_bnr_0')
// (12, 13, 'neigh_op_top_0')
// (12, 14, 'local_g3_0')
// (12, 14, 'lutff_0/in_1')
// (12, 14, 'lutff_0/out')
// (12, 15, 'neigh_op_bot_0')
// (13, 13, 'neigh_op_tnl_0')
// (13, 14, 'neigh_op_lft_0')
// (13, 15, 'neigh_op_bnl_0')

wire n443;
// (11, 13, 'neigh_op_tnr_1')
// (11, 14, 'neigh_op_rgt_1')
// (11, 15, 'neigh_op_bnr_1')
// (12, 13, 'neigh_op_top_1')
// (12, 14, 'local_g3_1')
// (12, 14, 'lutff_1/in_1')
// (12, 14, 'lutff_1/out')
// (12, 15, 'neigh_op_bot_1')
// (13, 13, 'neigh_op_tnl_1')
// (13, 14, 'neigh_op_lft_1')
// (13, 15, 'neigh_op_bnl_1')

wire n444;
// (11, 13, 'neigh_op_tnr_2')
// (11, 14, 'neigh_op_rgt_2')
// (11, 15, 'neigh_op_bnr_2')
// (12, 13, 'neigh_op_top_2')
// (12, 14, 'local_g3_2')
// (12, 14, 'lutff_2/in_1')
// (12, 14, 'lutff_2/out')
// (12, 15, 'neigh_op_bot_2')
// (13, 13, 'neigh_op_tnl_2')
// (13, 14, 'neigh_op_lft_2')
// (13, 15, 'neigh_op_bnl_2')

wire n445;
// (11, 13, 'neigh_op_tnr_3')
// (11, 14, 'neigh_op_rgt_3')
// (11, 14, 'sp4_r_v_b_38')
// (11, 15, 'neigh_op_bnr_3')
// (11, 15, 'sp4_r_v_b_27')
// (11, 16, 'sp4_r_v_b_14')
// (11, 17, 'sp4_r_v_b_3')
// (12, 13, 'neigh_op_top_3')
// (12, 13, 'sp4_v_t_38')
// (12, 14, 'local_g2_6')
// (12, 14, 'lutff_3/in_1')
// (12, 14, 'lutff_3/out')
// (12, 14, 'sp4_v_b_38')
// (12, 15, 'neigh_op_bot_3')
// (12, 15, 'sp4_v_b_27')
// (12, 16, 'sp4_v_b_14')
// (12, 17, 'sp4_v_b_3')
// (13, 13, 'neigh_op_tnl_3')
// (13, 14, 'neigh_op_lft_3')
// (13, 15, 'neigh_op_bnl_3')

wire n446;
// (11, 13, 'neigh_op_tnr_4')
// (11, 14, 'neigh_op_rgt_4')
// (11, 15, 'neigh_op_bnr_4')
// (12, 13, 'neigh_op_top_4')
// (12, 14, 'local_g3_4')
// (12, 14, 'lutff_4/in_1')
// (12, 14, 'lutff_4/out')
// (12, 15, 'neigh_op_bot_4')
// (13, 13, 'neigh_op_tnl_4')
// (13, 14, 'neigh_op_lft_4')
// (13, 15, 'neigh_op_bnl_4')

wire n447;
// (11, 13, 'neigh_op_tnr_5')
// (11, 14, 'neigh_op_rgt_5')
// (11, 15, 'neigh_op_bnr_5')
// (12, 13, 'neigh_op_top_5')
// (12, 14, 'local_g1_5')
// (12, 14, 'lutff_5/in_1')
// (12, 14, 'lutff_5/out')
// (12, 15, 'neigh_op_bot_5')
// (13, 13, 'neigh_op_tnl_5')
// (13, 14, 'neigh_op_lft_5')
// (13, 15, 'neigh_op_bnl_5')

wire n448;
// (11, 13, 'neigh_op_tnr_6')
// (11, 14, 'neigh_op_rgt_6')
// (11, 15, 'neigh_op_bnr_6')
// (12, 13, 'neigh_op_top_6')
// (12, 14, 'local_g1_6')
// (12, 14, 'lutff_6/in_1')
// (12, 14, 'lutff_6/out')
// (12, 15, 'neigh_op_bot_6')
// (13, 13, 'neigh_op_tnl_6')
// (13, 14, 'neigh_op_lft_6')
// (13, 15, 'neigh_op_bnl_6')

wire n449;
// (11, 13, 'neigh_op_tnr_7')
// (11, 14, 'neigh_op_rgt_7')
// (11, 15, 'neigh_op_bnr_7')
// (12, 13, 'neigh_op_top_7')
// (12, 14, 'local_g1_7')
// (12, 14, 'lutff_7/in_1')
// (12, 14, 'lutff_7/out')
// (12, 15, 'neigh_op_bot_7')
// (13, 13, 'neigh_op_tnl_7')
// (13, 14, 'neigh_op_lft_7')
// (13, 15, 'neigh_op_bnl_7')

reg n450 = 0;
// (11, 13, 'sp12_h_r_1')
// (12, 13, 'sp12_h_r_2')
// (13, 12, 'neigh_op_tnr_7')
// (13, 13, 'neigh_op_rgt_7')
// (13, 13, 'sp12_h_r_5')
// (13, 14, 'neigh_op_bnr_7')
// (14, 12, 'neigh_op_top_7')
// (14, 13, 'lutff_7/out')
// (14, 13, 'sp12_h_r_6')
// (14, 14, 'neigh_op_bot_7')
// (15, 12, 'neigh_op_tnl_7')
// (15, 13, 'neigh_op_lft_7')
// (15, 13, 'sp12_h_r_9')
// (15, 14, 'neigh_op_bnl_7')
// (16, 13, 'sp12_h_r_10')
// (17, 13, 'local_g1_5')
// (17, 13, 'lutff_7/in_3')
// (17, 13, 'sp12_h_r_13')
// (18, 13, 'sp12_h_r_14')
// (19, 13, 'sp12_h_r_17')
// (20, 13, 'sp12_h_r_18')
// (21, 13, 'sp12_h_r_21')
// (22, 13, 'sp12_h_r_22')
// (23, 13, 'sp12_h_l_22')

wire n451;
// (11, 14, 'lutff_0/cout')
// (11, 14, 'lutff_1/in_3')

wire n452;
// (11, 14, 'lutff_1/cout')
// (11, 14, 'lutff_2/in_3')

wire n453;
// (11, 14, 'lutff_2/cout')
// (11, 14, 'lutff_3/in_3')

wire n454;
// (11, 14, 'lutff_3/cout')
// (11, 14, 'lutff_4/in_3')

wire n455;
// (11, 14, 'lutff_4/cout')
// (11, 14, 'lutff_5/in_3')

wire n456;
// (11, 14, 'lutff_5/cout')
// (11, 14, 'lutff_6/in_3')

wire n457;
// (11, 14, 'lutff_6/cout')
// (11, 14, 'lutff_7/in_3')

wire n458;
// (11, 14, 'lutff_7/cout')
// (11, 15, 'carry_in')
// (11, 15, 'carry_in_mux')
// (11, 15, 'lutff_0/in_3')

wire n459;
// (11, 14, 'neigh_op_tnr_0')
// (11, 15, 'neigh_op_rgt_0')
// (11, 16, 'neigh_op_bnr_0')
// (12, 14, 'neigh_op_top_0')
// (12, 15, 'local_g3_0')
// (12, 15, 'lutff_0/in_1')
// (12, 15, 'lutff_0/out')
// (12, 16, 'neigh_op_bot_0')
// (13, 14, 'neigh_op_tnl_0')
// (13, 15, 'neigh_op_lft_0')
// (13, 16, 'neigh_op_bnl_0')

wire n460;
// (11, 14, 'neigh_op_tnr_1')
// (11, 15, 'neigh_op_rgt_1')
// (11, 16, 'neigh_op_bnr_1')
// (12, 14, 'neigh_op_top_1')
// (12, 15, 'local_g3_1')
// (12, 15, 'lutff_1/in_1')
// (12, 15, 'lutff_1/out')
// (12, 16, 'neigh_op_bot_1')
// (13, 14, 'neigh_op_tnl_1')
// (13, 15, 'neigh_op_lft_1')
// (13, 16, 'neigh_op_bnl_1')

wire n461;
// (11, 14, 'neigh_op_tnr_2')
// (11, 15, 'neigh_op_rgt_2')
// (11, 16, 'neigh_op_bnr_2')
// (12, 14, 'neigh_op_top_2')
// (12, 15, 'local_g3_2')
// (12, 15, 'lutff_2/in_1')
// (12, 15, 'lutff_2/out')
// (12, 16, 'neigh_op_bot_2')
// (13, 14, 'neigh_op_tnl_2')
// (13, 15, 'neigh_op_lft_2')
// (13, 16, 'neigh_op_bnl_2')

wire n462;
// (11, 14, 'neigh_op_tnr_3')
// (11, 15, 'neigh_op_rgt_3')
// (11, 16, 'neigh_op_bnr_3')
// (12, 14, 'neigh_op_top_3')
// (12, 15, 'local_g1_3')
// (12, 15, 'lutff_3/in_1')
// (12, 15, 'lutff_3/out')
// (12, 16, 'neigh_op_bot_3')
// (13, 14, 'neigh_op_tnl_3')
// (13, 15, 'neigh_op_lft_3')
// (13, 16, 'neigh_op_bnl_3')

wire n463;
// (11, 14, 'neigh_op_tnr_4')
// (11, 15, 'neigh_op_rgt_4')
// (11, 16, 'neigh_op_bnr_4')
// (12, 14, 'neigh_op_top_4')
// (12, 15, 'local_g1_4')
// (12, 15, 'lutff_4/in_1')
// (12, 15, 'lutff_4/out')
// (12, 16, 'neigh_op_bot_4')
// (13, 14, 'neigh_op_tnl_4')
// (13, 15, 'neigh_op_lft_4')
// (13, 16, 'neigh_op_bnl_4')

wire n464;
// (11, 14, 'neigh_op_tnr_5')
// (11, 15, 'neigh_op_rgt_5')
// (11, 16, 'neigh_op_bnr_5')
// (12, 14, 'neigh_op_top_5')
// (12, 15, 'local_g1_5')
// (12, 15, 'lutff_5/in_1')
// (12, 15, 'lutff_5/out')
// (12, 16, 'neigh_op_bot_5')
// (13, 14, 'neigh_op_tnl_5')
// (13, 15, 'neigh_op_lft_5')
// (13, 16, 'neigh_op_bnl_5')

wire n465;
// (11, 14, 'neigh_op_tnr_6')
// (11, 15, 'neigh_op_rgt_6')
// (11, 16, 'neigh_op_bnr_6')
// (12, 14, 'neigh_op_top_6')
// (12, 15, 'local_g1_6')
// (12, 15, 'lutff_6/in_1')
// (12, 15, 'lutff_6/out')
// (12, 16, 'neigh_op_bot_6')
// (13, 14, 'neigh_op_tnl_6')
// (13, 15, 'neigh_op_lft_6')
// (13, 16, 'neigh_op_bnl_6')

wire n466;
// (11, 14, 'neigh_op_tnr_7')
// (11, 15, 'neigh_op_rgt_7')
// (11, 16, 'neigh_op_bnr_7')
// (12, 14, 'neigh_op_top_7')
// (12, 15, 'local_g1_7')
// (12, 15, 'lutff_7/in_1')
// (12, 15, 'lutff_7/out')
// (12, 16, 'neigh_op_bot_7')
// (13, 14, 'neigh_op_tnl_7')
// (13, 15, 'neigh_op_lft_7')
// (13, 16, 'neigh_op_bnl_7')

wire n467;
// (11, 14, 'sp12_h_r_1')
// (12, 14, 'sp12_h_r_2')
// (13, 14, 'sp12_h_r_5')
// (14, 14, 'sp12_h_r_6')
// (15, 13, 'neigh_op_tnr_1')
// (15, 14, 'neigh_op_rgt_1')
// (15, 14, 'sp12_h_r_9')
// (15, 15, 'neigh_op_bnr_1')
// (16, 13, 'neigh_op_top_1')
// (16, 14, 'lutff_1/out')
// (16, 14, 'sp12_h_r_10')
// (16, 15, 'neigh_op_bot_1')
// (17, 13, 'neigh_op_tnl_1')
// (17, 14, 'neigh_op_lft_1')
// (17, 14, 'sp12_h_r_13')
// (17, 15, 'neigh_op_bnl_1')
// (18, 14, 'sp12_h_r_14')
// (19, 14, 'sp12_h_r_17')
// (20, 14, 'sp12_h_r_18')
// (21, 14, 'sp12_h_r_21')
// (22, 14, 'sp12_h_r_22')
// (23, 14, 'sp12_h_l_22')
// (23, 14, 'sp12_h_r_1')
// (24, 14, 'local_g0_2')
// (24, 14, 'lutff_global/cen')
// (24, 14, 'sp12_h_r_2')
// (25, 14, 'sp12_h_r_5')
// (26, 14, 'sp12_h_r_6')
// (27, 14, 'sp12_h_r_9')
// (28, 14, 'sp12_h_r_10')
// (29, 14, 'sp12_h_r_13')
// (30, 14, 'sp12_h_r_14')
// (31, 14, 'sp12_h_r_17')
// (32, 14, 'sp12_h_r_18')
// (33, 14, 'span12_horz_18')

reg n468 = 0;
// (11, 14, 'sp4_r_v_b_37')
// (11, 15, 'sp4_r_v_b_24')
// (11, 16, 'neigh_op_tnr_0')
// (11, 16, 'sp4_r_v_b_13')
// (11, 16, 'sp4_r_v_b_45')
// (11, 17, 'neigh_op_rgt_0')
// (11, 17, 'sp4_r_v_b_0')
// (11, 17, 'sp4_r_v_b_32')
// (11, 18, 'neigh_op_bnr_0')
// (11, 18, 'sp4_r_v_b_21')
// (11, 19, 'sp4_r_v_b_8')
// (12, 13, 'sp4_v_t_37')
// (12, 14, 'local_g2_5')
// (12, 14, 'lutff_0/in_3')
// (12, 14, 'sp4_v_b_37')
// (12, 15, 'sp4_v_b_24')
// (12, 15, 'sp4_v_t_45')
// (12, 16, 'neigh_op_top_0')
// (12, 16, 'sp4_v_b_13')
// (12, 16, 'sp4_v_b_45')
// (12, 17, 'local_g1_0')
// (12, 17, 'lutff_0/in_1')
// (12, 17, 'lutff_0/out')
// (12, 17, 'sp4_v_b_0')
// (12, 17, 'sp4_v_b_32')
// (12, 18, 'neigh_op_bot_0')
// (12, 18, 'sp4_v_b_21')
// (12, 19, 'sp4_h_r_8')
// (12, 19, 'sp4_v_b_8')
// (13, 16, 'neigh_op_tnl_0')
// (13, 17, 'neigh_op_lft_0')
// (13, 18, 'neigh_op_bnl_0')
// (13, 19, 'sp4_h_r_21')
// (14, 19, 'sp4_h_r_32')
// (15, 19, 'sp4_h_r_45')
// (15, 20, 'sp4_r_v_b_36')
// (15, 21, 'sp4_r_v_b_25')
// (15, 22, 'sp4_r_v_b_12')
// (15, 23, 'sp4_r_v_b_1')
// (16, 19, 'sp4_h_l_45')
// (16, 19, 'sp4_v_t_36')
// (16, 20, 'sp4_v_b_36')
// (16, 21, 'sp4_v_b_25')
// (16, 22, 'sp4_v_b_12')
// (16, 23, 'local_g1_1')
// (16, 23, 'lutff_5/in_3')
// (16, 23, 'sp4_v_b_1')

reg n469 = 0;
// (11, 14, 'sp4_r_v_b_39')
// (11, 15, 'sp4_r_v_b_26')
// (11, 16, 'neigh_op_tnr_1')
// (11, 16, 'sp4_r_v_b_15')
// (11, 16, 'sp4_r_v_b_47')
// (11, 17, 'neigh_op_rgt_1')
// (11, 17, 'sp4_r_v_b_2')
// (11, 17, 'sp4_r_v_b_34')
// (11, 18, 'neigh_op_bnr_1')
// (11, 18, 'sp4_r_v_b_23')
// (11, 19, 'sp4_r_v_b_10')
// (12, 13, 'sp4_v_t_39')
// (12, 14, 'local_g3_7')
// (12, 14, 'lutff_1/in_3')
// (12, 14, 'sp4_v_b_39')
// (12, 15, 'sp4_v_b_26')
// (12, 15, 'sp4_v_t_47')
// (12, 16, 'neigh_op_top_1')
// (12, 16, 'sp4_v_b_15')
// (12, 16, 'sp4_v_b_47')
// (12, 17, 'local_g3_1')
// (12, 17, 'lutff_1/in_1')
// (12, 17, 'lutff_1/out')
// (12, 17, 'sp4_v_b_2')
// (12, 17, 'sp4_v_b_34')
// (12, 18, 'neigh_op_bot_1')
// (12, 18, 'sp4_v_b_23')
// (12, 19, 'sp4_h_r_10')
// (12, 19, 'sp4_v_b_10')
// (13, 16, 'neigh_op_tnl_1')
// (13, 17, 'neigh_op_lft_1')
// (13, 18, 'neigh_op_bnl_1')
// (13, 19, 'sp4_h_r_23')
// (14, 19, 'sp4_h_r_34')
// (15, 19, 'sp4_h_r_47')
// (15, 20, 'sp4_r_v_b_47')
// (15, 21, 'sp4_r_v_b_34')
// (15, 22, 'sp4_r_v_b_23')
// (15, 23, 'sp4_r_v_b_10')
// (16, 19, 'sp4_h_l_47')
// (16, 19, 'sp4_v_t_47')
// (16, 20, 'sp4_v_b_47')
// (16, 21, 'sp4_v_b_34')
// (16, 22, 'sp4_v_b_23')
// (16, 23, 'local_g1_2')
// (16, 23, 'lutff_6/in_3')
// (16, 23, 'sp4_v_b_10')

reg n470 = 0;
// (11, 14, 'sp4_r_v_b_41')
// (11, 15, 'sp4_r_v_b_28')
// (11, 16, 'neigh_op_tnr_2')
// (11, 16, 'sp4_r_v_b_17')
// (11, 17, 'neigh_op_rgt_2')
// (11, 17, 'sp4_r_v_b_4')
// (11, 18, 'neigh_op_bnr_2')
// (12, 13, 'sp4_v_t_41')
// (12, 14, 'local_g2_1')
// (12, 14, 'lutff_2/in_3')
// (12, 14, 'sp4_v_b_41')
// (12, 15, 'sp4_v_b_28')
// (12, 16, 'neigh_op_top_2')
// (12, 16, 'sp4_v_b_17')
// (12, 17, 'local_g1_2')
// (12, 17, 'lutff_2/in_1')
// (12, 17, 'lutff_2/out')
// (12, 17, 'sp4_v_b_4')
// (12, 18, 'neigh_op_bot_2')
// (13, 16, 'neigh_op_tnl_2')
// (13, 17, 'neigh_op_lft_2')
// (13, 18, 'neigh_op_bnl_2')

reg n471 = 0;
// (11, 14, 'sp4_r_v_b_43')
// (11, 15, 'sp4_r_v_b_30')
// (11, 16, 'neigh_op_tnr_3')
// (11, 16, 'sp4_r_v_b_19')
// (11, 17, 'neigh_op_rgt_3')
// (11, 17, 'sp4_r_v_b_6')
// (11, 18, 'neigh_op_bnr_3')
// (12, 13, 'sp4_v_t_43')
// (12, 14, 'local_g3_3')
// (12, 14, 'lutff_3/in_3')
// (12, 14, 'sp4_v_b_43')
// (12, 15, 'sp4_v_b_30')
// (12, 16, 'neigh_op_top_3')
// (12, 16, 'sp4_v_b_19')
// (12, 17, 'local_g1_3')
// (12, 17, 'lutff_3/in_1')
// (12, 17, 'lutff_3/out')
// (12, 17, 'sp4_v_b_6')
// (12, 18, 'neigh_op_bot_3')
// (13, 16, 'neigh_op_tnl_3')
// (13, 17, 'neigh_op_lft_3')
// (13, 18, 'neigh_op_bnl_3')

reg n472 = 0;
// (11, 14, 'sp4_r_v_b_45')
// (11, 15, 'sp4_r_v_b_32')
// (11, 16, 'neigh_op_tnr_4')
// (11, 16, 'sp4_r_v_b_21')
// (11, 17, 'neigh_op_rgt_4')
// (11, 17, 'sp4_r_v_b_8')
// (11, 18, 'neigh_op_bnr_4')
// (12, 13, 'sp4_v_t_45')
// (12, 14, 'local_g3_5')
// (12, 14, 'lutff_4/in_0')
// (12, 14, 'sp4_v_b_45')
// (12, 15, 'sp4_v_b_32')
// (12, 16, 'neigh_op_top_4')
// (12, 16, 'sp4_v_b_21')
// (12, 17, 'local_g3_4')
// (12, 17, 'lutff_4/in_1')
// (12, 17, 'lutff_4/out')
// (12, 17, 'sp4_v_b_8')
// (12, 18, 'neigh_op_bot_4')
// (13, 16, 'neigh_op_tnl_4')
// (13, 17, 'neigh_op_lft_4')
// (13, 18, 'neigh_op_bnl_4')

reg n473 = 0;
// (11, 14, 'sp4_r_v_b_47')
// (11, 15, 'sp4_r_v_b_34')
// (11, 16, 'neigh_op_tnr_5')
// (11, 16, 'sp4_r_v_b_23')
// (11, 17, 'neigh_op_rgt_5')
// (11, 17, 'sp4_r_v_b_10')
// (11, 18, 'neigh_op_bnr_5')
// (12, 13, 'sp4_v_t_47')
// (12, 14, 'local_g2_7')
// (12, 14, 'lutff_5/in_0')
// (12, 14, 'sp4_v_b_47')
// (12, 15, 'sp4_v_b_34')
// (12, 16, 'neigh_op_top_5')
// (12, 16, 'sp4_v_b_23')
// (12, 17, 'local_g3_5')
// (12, 17, 'lutff_5/in_1')
// (12, 17, 'lutff_5/out')
// (12, 17, 'sp4_v_b_10')
// (12, 18, 'neigh_op_bot_5')
// (13, 16, 'neigh_op_tnl_5')
// (13, 17, 'neigh_op_lft_5')
// (13, 18, 'neigh_op_bnl_5')

wire n474;
// (11, 15, 'lutff_0/cout')
// (11, 15, 'lutff_1/in_3')

wire n475;
// (11, 15, 'lutff_1/cout')
// (11, 15, 'lutff_2/in_3')

wire n476;
// (11, 15, 'lutff_2/cout')
// (11, 15, 'lutff_3/in_3')

wire n477;
// (11, 15, 'lutff_3/cout')
// (11, 15, 'lutff_4/in_3')

wire n478;
// (11, 15, 'lutff_4/cout')
// (11, 15, 'lutff_5/in_3')

wire n479;
// (11, 15, 'lutff_5/cout')
// (11, 15, 'lutff_6/in_3')

wire n480;
// (11, 15, 'lutff_6/cout')
// (11, 15, 'lutff_7/in_3')

wire n481;
// (11, 15, 'neigh_op_tnr_0')
// (11, 16, 'local_g3_0')
// (11, 16, 'lutff_0/in_3')
// (11, 16, 'neigh_op_rgt_0')
// (11, 17, 'neigh_op_bnr_0')
// (12, 15, 'neigh_op_top_0')
// (12, 16, 'local_g2_0')
// (12, 16, 'lutff_0/out')
// (12, 16, 'lutff_5/in_3')
// (12, 17, 'neigh_op_bot_0')
// (13, 15, 'neigh_op_tnl_0')
// (13, 16, 'neigh_op_lft_0')
// (13, 17, 'neigh_op_bnl_0')

wire n482;
// (11, 15, 'neigh_op_tnr_5')
// (11, 16, 'neigh_op_rgt_5')
// (11, 17, 'local_g1_5')
// (11, 17, 'lutff_5/in_3')
// (11, 17, 'neigh_op_bnr_5')
// (12, 15, 'neigh_op_top_5')
// (12, 16, 'lutff_5/out')
// (12, 17, 'neigh_op_bot_5')
// (13, 15, 'neigh_op_tnl_5')
// (13, 16, 'neigh_op_lft_5')
// (13, 17, 'neigh_op_bnl_5')

reg n483 = 0;
// (11, 15, 'sp12_h_r_0')
// (12, 15, 'sp12_h_r_3')
// (13, 15, 'sp12_h_r_4')
// (14, 14, 'neigh_op_tnr_0')
// (14, 15, 'neigh_op_rgt_0')
// (14, 15, 'sp12_h_r_7')
// (14, 16, 'neigh_op_bnr_0')
// (15, 14, 'neigh_op_top_0')
// (15, 15, 'lutff_0/out')
// (15, 15, 'sp12_h_r_8')
// (15, 16, 'neigh_op_bot_0')
// (16, 14, 'neigh_op_tnl_0')
// (16, 15, 'neigh_op_lft_0')
// (16, 15, 'sp12_h_r_11')
// (16, 16, 'neigh_op_bnl_0')
// (17, 15, 'sp12_h_r_12')
// (18, 15, 'local_g1_7')
// (18, 15, 'lutff_3/in_1')
// (18, 15, 'sp12_h_r_15')
// (19, 15, 'sp12_h_r_16')
// (20, 15, 'sp12_h_r_19')
// (21, 15, 'sp12_h_r_20')
// (22, 15, 'sp12_h_r_23')
// (23, 15, 'sp12_h_l_23')

reg n484 = 0;
// (11, 15, 'sp4_r_v_b_37')
// (11, 16, 'sp4_r_v_b_24')
// (11, 17, 'neigh_op_tnr_0')
// (11, 17, 'sp4_r_v_b_13')
// (11, 18, 'neigh_op_rgt_0')
// (11, 18, 'sp4_r_v_b_0')
// (11, 19, 'neigh_op_bnr_0')
// (12, 14, 'sp4_v_t_37')
// (12, 15, 'local_g2_5')
// (12, 15, 'lutff_0/in_3')
// (12, 15, 'sp4_v_b_37')
// (12, 16, 'sp4_v_b_24')
// (12, 17, 'neigh_op_top_0')
// (12, 17, 'sp4_v_b_13')
// (12, 18, 'local_g3_0')
// (12, 18, 'lutff_0/in_1')
// (12, 18, 'lutff_0/out')
// (12, 18, 'sp4_v_b_0')
// (12, 19, 'neigh_op_bot_0')
// (13, 17, 'neigh_op_tnl_0')
// (13, 18, 'neigh_op_lft_0')
// (13, 19, 'neigh_op_bnl_0')

reg n485 = 0;
// (11, 15, 'sp4_r_v_b_39')
// (11, 16, 'sp4_r_v_b_26')
// (11, 17, 'neigh_op_tnr_1')
// (11, 17, 'sp4_r_v_b_15')
// (11, 18, 'neigh_op_rgt_1')
// (11, 18, 'sp4_r_v_b_2')
// (11, 19, 'neigh_op_bnr_1')
// (12, 14, 'sp4_v_t_39')
// (12, 15, 'local_g3_7')
// (12, 15, 'lutff_1/in_3')
// (12, 15, 'sp4_v_b_39')
// (12, 16, 'sp4_v_b_26')
// (12, 17, 'neigh_op_top_1')
// (12, 17, 'sp4_v_b_15')
// (12, 18, 'local_g3_1')
// (12, 18, 'lutff_1/in_1')
// (12, 18, 'lutff_1/out')
// (12, 18, 'sp4_v_b_2')
// (12, 19, 'neigh_op_bot_1')
// (13, 17, 'neigh_op_tnl_1')
// (13, 18, 'neigh_op_lft_1')
// (13, 19, 'neigh_op_bnl_1')

reg n486 = 0;
// (11, 15, 'sp4_r_v_b_41')
// (11, 16, 'sp4_r_v_b_28')
// (11, 17, 'neigh_op_tnr_2')
// (11, 17, 'sp4_r_v_b_17')
// (11, 18, 'neigh_op_rgt_2')
// (11, 18, 'sp4_r_v_b_4')
// (11, 19, 'neigh_op_bnr_2')
// (12, 14, 'sp4_v_t_41')
// (12, 15, 'local_g2_1')
// (12, 15, 'lutff_2/in_3')
// (12, 15, 'sp4_v_b_41')
// (12, 16, 'sp4_v_b_28')
// (12, 17, 'neigh_op_top_2')
// (12, 17, 'sp4_v_b_17')
// (12, 18, 'local_g1_2')
// (12, 18, 'lutff_2/in_1')
// (12, 18, 'lutff_2/out')
// (12, 18, 'sp4_v_b_4')
// (12, 19, 'neigh_op_bot_2')
// (13, 17, 'neigh_op_tnl_2')
// (13, 18, 'neigh_op_lft_2')
// (13, 19, 'neigh_op_bnl_2')

reg n487 = 0;
// (11, 15, 'sp4_r_v_b_43')
// (11, 16, 'sp4_r_v_b_30')
// (11, 17, 'neigh_op_tnr_3')
// (11, 17, 'sp4_r_v_b_19')
// (11, 18, 'neigh_op_rgt_3')
// (11, 18, 'sp4_r_v_b_6')
// (11, 19, 'neigh_op_bnr_3')
// (12, 14, 'sp4_v_t_43')
// (12, 15, 'local_g3_3')
// (12, 15, 'lutff_3/in_3')
// (12, 15, 'sp4_v_b_43')
// (12, 16, 'sp4_v_b_30')
// (12, 17, 'neigh_op_top_3')
// (12, 17, 'sp4_v_b_19')
// (12, 18, 'local_g1_3')
// (12, 18, 'lutff_3/in_1')
// (12, 18, 'lutff_3/out')
// (12, 18, 'sp4_v_b_6')
// (12, 19, 'neigh_op_bot_3')
// (13, 17, 'neigh_op_tnl_3')
// (13, 18, 'neigh_op_lft_3')
// (13, 19, 'neigh_op_bnl_3')

reg n488 = 0;
// (11, 15, 'sp4_r_v_b_47')
// (11, 16, 'sp4_r_v_b_34')
// (11, 17, 'neigh_op_tnr_5')
// (11, 17, 'sp4_r_v_b_23')
// (11, 18, 'neigh_op_rgt_5')
// (11, 18, 'sp4_r_v_b_10')
// (11, 19, 'neigh_op_bnr_5')
// (12, 14, 'sp4_v_t_47')
// (12, 15, 'local_g2_7')
// (12, 15, 'lutff_5/in_0')
// (12, 15, 'sp4_v_b_47')
// (12, 16, 'sp4_v_b_34')
// (12, 17, 'neigh_op_top_5')
// (12, 17, 'sp4_v_b_23')
// (12, 18, 'local_g1_5')
// (12, 18, 'lutff_5/in_1')
// (12, 18, 'lutff_5/out')
// (12, 18, 'sp4_v_b_10')
// (12, 19, 'neigh_op_bot_5')
// (13, 17, 'neigh_op_tnl_5')
// (13, 18, 'neigh_op_lft_5')
// (13, 19, 'neigh_op_bnl_5')

wire n489;
// (11, 16, 'lutff_0/lout')
// (11, 16, 'lutff_1/in_2')

reg n490 = 0;
// (11, 16, 'neigh_op_tnr_6')
// (11, 17, 'neigh_op_rgt_6')
// (11, 18, 'neigh_op_bnr_6')
// (12, 11, 'sp12_v_t_23')
// (12, 12, 'sp12_v_b_23')
// (12, 13, 'sp12_v_b_20')
// (12, 14, 'local_g2_3')
// (12, 14, 'lutff_6/in_3')
// (12, 14, 'sp12_v_b_19')
// (12, 15, 'sp12_v_b_16')
// (12, 16, 'neigh_op_top_6')
// (12, 16, 'sp12_v_b_15')
// (12, 17, 'local_g1_6')
// (12, 17, 'lutff_6/in_1')
// (12, 17, 'lutff_6/out')
// (12, 17, 'sp12_v_b_12')
// (12, 18, 'neigh_op_bot_6')
// (12, 18, 'sp12_v_b_11')
// (12, 19, 'sp12_v_b_8')
// (12, 20, 'sp12_v_b_7')
// (12, 21, 'sp12_v_b_4')
// (12, 22, 'sp12_v_b_3')
// (12, 23, 'sp12_v_b_0')
// (13, 16, 'neigh_op_tnl_6')
// (13, 17, 'neigh_op_lft_6')
// (13, 18, 'neigh_op_bnl_6')

reg n491 = 0;
// (11, 16, 'neigh_op_tnr_7')
// (11, 17, 'neigh_op_rgt_7')
// (11, 18, 'neigh_op_bnr_7')
// (12, 13, 'sp4_r_v_b_47')
// (12, 14, 'local_g2_2')
// (12, 14, 'lutff_7/in_3')
// (12, 14, 'sp4_r_v_b_34')
// (12, 15, 'sp4_r_v_b_23')
// (12, 16, 'neigh_op_top_7')
// (12, 16, 'sp4_r_v_b_10')
// (12, 17, 'local_g3_7')
// (12, 17, 'lutff_7/in_1')
// (12, 17, 'lutff_7/out')
// (12, 17, 'sp4_r_v_b_47')
// (12, 18, 'neigh_op_bot_7')
// (12, 18, 'sp4_r_v_b_34')
// (12, 19, 'sp4_r_v_b_23')
// (12, 20, 'sp4_r_v_b_10')
// (13, 12, 'sp4_v_t_47')
// (13, 13, 'sp4_v_b_47')
// (13, 14, 'sp4_v_b_34')
// (13, 15, 'sp4_v_b_23')
// (13, 16, 'neigh_op_tnl_7')
// (13, 16, 'sp4_v_b_10')
// (13, 16, 'sp4_v_t_47')
// (13, 17, 'neigh_op_lft_7')
// (13, 17, 'sp4_v_b_47')
// (13, 18, 'neigh_op_bnl_7')
// (13, 18, 'sp4_v_b_34')
// (13, 19, 'sp4_v_b_23')
// (13, 20, 'sp4_v_b_10')

wire n492;
// (11, 16, 'sp4_h_r_11')
// (12, 16, 'sp4_h_r_22')
// (13, 16, 'local_g3_3')
// (13, 16, 'lutff_global/cen')
// (13, 16, 'sp4_h_r_35')
// (14, 15, 'neigh_op_tnr_4')
// (14, 16, 'neigh_op_rgt_4')
// (14, 16, 'sp4_h_r_46')
// (14, 17, 'neigh_op_bnr_4')
// (15, 15, 'neigh_op_top_4')
// (15, 16, 'lutff_4/out')
// (15, 16, 'sp4_h_l_46')
// (15, 16, 'sp4_h_r_8')
// (15, 17, 'neigh_op_bot_4')
// (16, 15, 'neigh_op_tnl_4')
// (16, 16, 'neigh_op_lft_4')
// (16, 16, 'sp4_h_r_21')
// (16, 17, 'neigh_op_bnl_4')
// (17, 16, 'sp4_h_r_32')
// (18, 16, 'sp4_h_r_45')
// (19, 16, 'sp4_h_l_45')

wire n493;
// (11, 17, 'local_g0_0')
// (11, 17, 'lutff_5/in_1')
// (11, 17, 'sp4_h_r_0')
// (12, 16, 'neigh_op_tnr_4')
// (12, 17, 'neigh_op_rgt_4')
// (12, 17, 'sp4_h_r_13')
// (12, 18, 'neigh_op_bnr_4')
// (13, 16, 'neigh_op_top_4')
// (13, 17, 'lutff_4/out')
// (13, 17, 'sp4_h_r_24')
// (13, 18, 'neigh_op_bot_4')
// (14, 16, 'neigh_op_tnl_4')
// (14, 17, 'neigh_op_lft_4')
// (14, 17, 'sp4_h_r_37')
// (14, 18, 'neigh_op_bnl_4')
// (15, 17, 'sp4_h_l_37')

reg n494 = 0;
// (11, 17, 'local_g0_2')
// (11, 17, 'lutff_3/in_3')
// (11, 17, 'sp4_h_r_2')
// (11, 18, 'local_g0_3')
// (11, 18, 'lutff_3/in_2')
// (11, 18, 'sp4_h_r_3')
// (11, 21, 'sp4_h_r_7')
// (12, 17, 'sp4_h_r_15')
// (12, 18, 'sp4_h_r_14')
// (12, 19, 'sp4_r_v_b_40')
// (12, 20, 'sp4_r_v_b_29')
// (12, 21, 'local_g0_2')
// (12, 21, 'lutff_3/in_1')
// (12, 21, 'sp4_h_r_18')
// (12, 21, 'sp4_r_v_b_16')
// (12, 22, 'sp4_r_v_b_5')
// (13, 17, 'local_g3_3')
// (13, 17, 'lutff_0/in_0')
// (13, 17, 'lutff_1/in_3')
// (13, 17, 'neigh_op_tnr_3')
// (13, 17, 'sp4_h_r_26')
// (13, 18, 'local_g3_3')
// (13, 18, 'lutff_3/in_3')
// (13, 18, 'neigh_op_rgt_3')
// (13, 18, 'sp4_h_r_11')
// (13, 18, 'sp4_h_r_27')
// (13, 18, 'sp4_v_t_40')
// (13, 19, 'neigh_op_bnr_3')
// (13, 19, 'sp4_v_b_40')
// (13, 20, 'sp4_v_b_29')
// (13, 21, 'sp4_h_r_31')
// (13, 21, 'sp4_v_b_16')
// (13, 22, 'local_g0_5')
// (13, 22, 'lutff_3/in_2')
// (13, 22, 'sp4_v_b_5')
// (14, 17, 'neigh_op_top_3')
// (14, 17, 'sp4_h_r_39')
// (14, 18, 'local_g1_3')
// (14, 18, 'lutff_3/in_1')
// (14, 18, 'lutff_3/out')
// (14, 18, 'sp4_h_r_22')
// (14, 18, 'sp4_h_r_38')
// (14, 18, 'sp4_r_v_b_39')
// (14, 19, 'neigh_op_bot_3')
// (14, 19, 'sp4_r_v_b_26')
// (14, 20, 'sp4_r_v_b_15')
// (14, 21, 'sp4_h_r_42')
// (14, 21, 'sp4_r_v_b_2')
// (15, 17, 'neigh_op_tnl_3')
// (15, 17, 'sp4_h_l_39')
// (15, 17, 'sp4_v_t_39')
// (15, 18, 'neigh_op_lft_3')
// (15, 18, 'sp4_h_l_38')
// (15, 18, 'sp4_h_r_35')
// (15, 18, 'sp4_v_b_39')
// (15, 19, 'neigh_op_bnl_3')
// (15, 19, 'sp4_v_b_26')
// (15, 20, 'local_g0_7')
// (15, 20, 'lutff_3/in_2')
// (15, 20, 'sp4_v_b_15')
// (15, 21, 'sp4_h_l_42')
// (15, 21, 'sp4_v_b_2')
// (16, 18, 'sp4_h_r_46')
// (16, 19, 'sp4_r_v_b_46')
// (16, 20, 'sp4_r_v_b_35')
// (16, 21, 'sp4_r_v_b_22')
// (16, 22, 'sp4_r_v_b_11')
// (17, 18, 'sp4_h_l_46')
// (17, 18, 'sp4_v_t_46')
// (17, 19, 'sp4_v_b_46')
// (17, 20, 'sp4_v_b_35')
// (17, 21, 'sp4_v_b_22')
// (17, 22, 'local_g1_3')
// (17, 22, 'lutff_3/in_1')
// (17, 22, 'sp4_v_b_11')

wire n495;
// (11, 17, 'local_g0_4')
// (11, 17, 'lutff_3/in_1')
// (11, 17, 'lutff_7/in_3')
// (11, 17, 'sp4_h_r_4')
// (12, 16, 'neigh_op_tnr_6')
// (12, 17, 'neigh_op_rgt_6')
// (12, 17, 'sp4_h_r_17')
// (12, 18, 'neigh_op_bnr_6')
// (13, 11, 'sp12_v_t_23')
// (13, 12, 'sp12_v_b_23')
// (13, 13, 'sp12_v_b_20')
// (13, 14, 'sp12_v_b_19')
// (13, 15, 'sp12_v_b_16')
// (13, 16, 'neigh_op_top_6')
// (13, 16, 'sp12_v_b_15')
// (13, 17, 'lutff_6/out')
// (13, 17, 'sp12_v_b_12')
// (13, 17, 'sp4_h_r_28')
// (13, 18, 'neigh_op_bot_6')
// (13, 18, 'sp12_v_b_11')
// (13, 19, 'sp12_v_b_8')
// (13, 20, 'sp12_v_b_7')
// (13, 21, 'local_g3_4')
// (13, 21, 'lutff_3/in_0')
// (13, 21, 'sp12_v_b_4')
// (13, 22, 'sp12_v_b_3')
// (13, 23, 'sp12_v_b_0')
// (14, 16, 'neigh_op_tnl_6')
// (14, 17, 'neigh_op_lft_6')
// (14, 17, 'sp4_h_r_41')
// (14, 18, 'neigh_op_bnl_6')
// (15, 17, 'sp4_h_l_41')

wire n496;
// (11, 17, 'lutff_3/lout')
// (11, 17, 'lutff_4/in_2')

wire n497;
// (11, 17, 'lutff_4/lout')
// (11, 17, 'lutff_5/in_2')

wire n498;
// (11, 17, 'lutff_6/lout')
// (11, 17, 'lutff_7/in_2')

reg n499 = 0;
// (11, 17, 'neigh_op_tnr_4')
// (11, 18, 'neigh_op_rgt_4')
// (11, 19, 'neigh_op_bnr_4')
// (12, 15, 'local_g3_4')
// (12, 15, 'lutff_4/in_3')
// (12, 15, 'sp4_r_v_b_44')
// (12, 16, 'sp4_r_v_b_33')
// (12, 17, 'neigh_op_top_4')
// (12, 17, 'sp4_r_v_b_20')
// (12, 18, 'local_g3_4')
// (12, 18, 'lutff_4/in_1')
// (12, 18, 'lutff_4/out')
// (12, 18, 'sp4_r_v_b_9')
// (12, 19, 'neigh_op_bot_4')
// (13, 14, 'sp4_v_t_44')
// (13, 15, 'sp4_v_b_44')
// (13, 16, 'sp4_v_b_33')
// (13, 17, 'neigh_op_tnl_4')
// (13, 17, 'sp4_v_b_20')
// (13, 18, 'neigh_op_lft_4')
// (13, 18, 'sp4_v_b_9')
// (13, 19, 'neigh_op_bnl_4')

reg n500 = 0;
// (11, 17, 'neigh_op_tnr_6')
// (11, 18, 'neigh_op_rgt_6')
// (11, 19, 'neigh_op_bnr_6')
// (12, 12, 'sp12_v_t_23')
// (12, 13, 'sp12_v_b_23')
// (12, 14, 'sp12_v_b_20')
// (12, 15, 'local_g2_3')
// (12, 15, 'lutff_6/in_3')
// (12, 15, 'sp12_v_b_19')
// (12, 16, 'sp12_v_b_16')
// (12, 17, 'neigh_op_top_6')
// (12, 17, 'sp12_v_b_15')
// (12, 18, 'local_g1_6')
// (12, 18, 'lutff_6/in_1')
// (12, 18, 'lutff_6/out')
// (12, 18, 'sp12_v_b_12')
// (12, 19, 'neigh_op_bot_6')
// (12, 19, 'sp12_v_b_11')
// (12, 20, 'sp12_v_b_8')
// (12, 21, 'sp12_v_b_7')
// (12, 22, 'sp12_v_b_4')
// (12, 23, 'sp12_v_b_3')
// (12, 24, 'sp12_v_b_0')
// (13, 17, 'neigh_op_tnl_6')
// (13, 18, 'neigh_op_lft_6')
// (13, 19, 'neigh_op_bnl_6')

reg n501 = 0;
// (11, 17, 'neigh_op_tnr_7')
// (11, 18, 'neigh_op_rgt_7')
// (11, 19, 'neigh_op_bnr_7')
// (12, 13, 'sp12_v_t_22')
// (12, 14, 'sp12_v_b_22')
// (12, 15, 'local_g3_5')
// (12, 15, 'lutff_7/in_3')
// (12, 15, 'sp12_v_b_21')
// (12, 16, 'sp12_v_b_18')
// (12, 17, 'neigh_op_top_7')
// (12, 17, 'sp12_v_b_17')
// (12, 18, 'local_g1_7')
// (12, 18, 'lutff_7/in_1')
// (12, 18, 'lutff_7/out')
// (12, 18, 'sp12_v_b_14')
// (12, 19, 'neigh_op_bot_7')
// (12, 19, 'sp12_v_b_13')
// (12, 20, 'sp12_v_b_10')
// (12, 21, 'sp12_v_b_9')
// (12, 22, 'sp12_v_b_6')
// (12, 23, 'sp12_v_b_5')
// (12, 24, 'sp12_v_b_2')
// (12, 25, 'sp12_v_b_1')
// (13, 17, 'neigh_op_tnl_7')
// (13, 18, 'neigh_op_lft_7')
// (13, 19, 'neigh_op_bnl_7')

reg n502 = 0;
// (11, 17, 'sp12_h_r_1')
// (12, 17, 'sp12_h_r_2')
// (13, 17, 'sp12_h_r_5')
// (14, 17, 'sp12_h_r_6')
// (15, 17, 'sp12_h_r_9')
// (16, 17, 'sp12_h_r_10')
// (17, 17, 'sp12_h_r_13')
// (18, 17, 'sp12_h_r_14')
// (19, 17, 'local_g0_1')
// (19, 17, 'lutff_2/in_1')
// (19, 17, 'sp12_h_r_17')
// (20, 17, 'sp12_h_r_18')
// (21, 17, 'sp12_h_r_21')
// (22, 11, 'neigh_op_tnr_5')
// (22, 12, 'neigh_op_rgt_5')
// (22, 13, 'neigh_op_bnr_5')
// (22, 17, 'sp12_h_r_22')
// (23, 5, 'sp12_v_t_22')
// (23, 6, 'sp12_v_b_22')
// (23, 7, 'sp12_v_b_21')
// (23, 8, 'sp12_v_b_18')
// (23, 9, 'sp12_v_b_17')
// (23, 10, 'sp12_v_b_14')
// (23, 11, 'neigh_op_top_5')
// (23, 11, 'sp12_v_b_13')
// (23, 12, 'lutff_5/out')
// (23, 12, 'sp12_v_b_10')
// (23, 13, 'neigh_op_bot_5')
// (23, 13, 'sp12_v_b_9')
// (23, 14, 'sp12_v_b_6')
// (23, 15, 'sp12_v_b_5')
// (23, 16, 'sp12_v_b_2')
// (23, 17, 'sp12_h_l_22')
// (23, 17, 'sp12_v_b_1')
// (24, 11, 'neigh_op_tnl_5')
// (24, 12, 'neigh_op_lft_5')
// (24, 13, 'neigh_op_bnl_5')

reg n503 = 0;
// (11, 18, 'local_g2_0')
// (11, 18, 'lutff_0/in_0')
// (11, 18, 'neigh_op_tnr_0')
// (11, 19, 'neigh_op_rgt_0')
// (11, 20, 'neigh_op_bnr_0')
// (12, 18, 'neigh_op_top_0')
// (12, 19, 'lutff_0/out')
// (12, 20, 'neigh_op_bot_0')
// (13, 18, 'neigh_op_tnl_0')
// (13, 19, 'neigh_op_lft_0')
// (13, 20, 'neigh_op_bnl_0')

reg n504 = 0;
// (11, 18, 'local_g3_1')
// (11, 18, 'lutff_1/in_3')
// (11, 18, 'neigh_op_tnr_1')
// (11, 19, 'neigh_op_rgt_1')
// (11, 20, 'neigh_op_bnr_1')
// (12, 18, 'neigh_op_top_1')
// (12, 19, 'lutff_1/out')
// (12, 20, 'neigh_op_bot_1')
// (13, 18, 'neigh_op_tnl_1')
// (13, 19, 'neigh_op_lft_1')
// (13, 20, 'neigh_op_bnl_1')

reg n505 = 0;
// (11, 18, 'local_g3_2')
// (11, 18, 'lutff_2/in_3')
// (11, 18, 'neigh_op_tnr_2')
// (11, 19, 'neigh_op_rgt_2')
// (11, 20, 'neigh_op_bnr_2')
// (12, 18, 'neigh_op_top_2')
// (12, 19, 'lutff_2/out')
// (12, 20, 'neigh_op_bot_2')
// (13, 18, 'neigh_op_tnl_2')
// (13, 19, 'neigh_op_lft_2')
// (13, 20, 'neigh_op_bnl_2')

reg n506 = 0;
// (11, 18, 'local_g3_3')
// (11, 18, 'lutff_3/in_3')
// (11, 18, 'neigh_op_tnr_3')
// (11, 19, 'neigh_op_rgt_3')
// (11, 20, 'neigh_op_bnr_3')
// (12, 18, 'neigh_op_top_3')
// (12, 19, 'lutff_3/out')
// (12, 20, 'neigh_op_bot_3')
// (13, 18, 'neigh_op_tnl_3')
// (13, 19, 'neigh_op_lft_3')
// (13, 20, 'neigh_op_bnl_3')

reg n507 = 0;
// (11, 18, 'local_g3_4')
// (11, 18, 'lutff_4/in_3')
// (11, 18, 'neigh_op_tnr_4')
// (11, 19, 'neigh_op_rgt_4')
// (11, 20, 'neigh_op_bnr_4')
// (12, 18, 'neigh_op_top_4')
// (12, 19, 'lutff_4/out')
// (12, 20, 'neigh_op_bot_4')
// (13, 18, 'neigh_op_tnl_4')
// (13, 19, 'neigh_op_lft_4')
// (13, 20, 'neigh_op_bnl_4')

reg n508 = 0;
// (11, 18, 'local_g3_5')
// (11, 18, 'lutff_5/in_3')
// (11, 18, 'neigh_op_tnr_5')
// (11, 19, 'neigh_op_rgt_5')
// (11, 20, 'neigh_op_bnr_5')
// (12, 18, 'neigh_op_top_5')
// (12, 19, 'lutff_5/out')
// (12, 20, 'neigh_op_bot_5')
// (13, 18, 'neigh_op_tnl_5')
// (13, 19, 'neigh_op_lft_5')
// (13, 20, 'neigh_op_bnl_5')

reg n509 = 0;
// (11, 18, 'local_g3_6')
// (11, 18, 'lutff_6/in_3')
// (11, 18, 'neigh_op_tnr_6')
// (11, 19, 'neigh_op_rgt_6')
// (11, 20, 'neigh_op_bnr_6')
// (12, 18, 'neigh_op_top_6')
// (12, 19, 'lutff_6/out')
// (12, 20, 'neigh_op_bot_6')
// (13, 18, 'neigh_op_tnl_6')
// (13, 19, 'neigh_op_lft_6')
// (13, 20, 'neigh_op_bnl_6')

reg n510 = 0;
// (11, 18, 'local_g3_7')
// (11, 18, 'lutff_7/in_3')
// (11, 18, 'neigh_op_tnr_7')
// (11, 19, 'neigh_op_rgt_7')
// (11, 20, 'neigh_op_bnr_7')
// (12, 18, 'neigh_op_top_7')
// (12, 19, 'lutff_7/out')
// (12, 20, 'neigh_op_bot_7')
// (13, 18, 'neigh_op_tnl_7')
// (13, 19, 'neigh_op_lft_7')
// (13, 20, 'neigh_op_bnl_7')

wire n511;
// (11, 18, 'lutff_7/cout')
// (11, 19, 'carry_in')
// (11, 19, 'carry_in_mux')

wire n512;
// (11, 18, 'sp12_h_r_0')
// (12, 17, 'neigh_op_tnr_6')
// (12, 18, 'neigh_op_rgt_6')
// (12, 18, 'sp12_h_r_3')
// (12, 19, 'neigh_op_bnr_6')
// (13, 17, 'neigh_op_top_6')
// (13, 18, 'local_g2_6')
// (13, 18, 'lutff_6/in_2')
// (13, 18, 'lutff_6/out')
// (13, 18, 'sp12_h_r_4')
// (13, 19, 'neigh_op_bot_6')
// (14, 17, 'neigh_op_tnl_6')
// (14, 18, 'neigh_op_lft_6')
// (14, 18, 'sp12_h_r_7')
// (14, 19, 'neigh_op_bnl_6')
// (15, 18, 'sp12_h_r_8')
// (16, 18, 'sp12_h_r_11')
// (17, 18, 'local_g0_4')
// (17, 18, 'lutff_6/in_2')
// (17, 18, 'sp12_h_r_12')
// (18, 18, 'sp12_h_r_15')
// (19, 18, 'sp12_h_r_16')
// (20, 18, 'sp12_h_r_19')
// (21, 18, 'sp12_h_r_20')
// (22, 18, 'sp12_h_r_23')
// (23, 18, 'sp12_h_l_23')

reg n513 = 0;
// (11, 19, 'local_g0_1')
// (11, 19, 'lutff_7/in_2')
// (11, 19, 'sp12_h_r_1')
// (12, 19, 'sp12_h_r_2')
// (12, 20, 'sp4_r_v_b_38')
// (12, 21, 'sp4_r_v_b_27')
// (12, 22, 'local_g2_6')
// (12, 22, 'lutff_7/in_1')
// (12, 22, 'sp4_r_v_b_14')
// (12, 23, 'sp4_r_v_b_3')
// (13, 17, 'sp4_r_v_b_38')
// (13, 18, 'neigh_op_tnr_7')
// (13, 18, 'sp4_r_v_b_27')
// (13, 18, 'sp4_r_v_b_43')
// (13, 19, 'local_g3_7')
// (13, 19, 'lutff_7/in_3')
// (13, 19, 'neigh_op_rgt_7')
// (13, 19, 'sp12_h_r_5')
// (13, 19, 'sp4_h_r_3')
// (13, 19, 'sp4_r_v_b_14')
// (13, 19, 'sp4_r_v_b_30')
// (13, 19, 'sp4_v_t_38')
// (13, 20, 'neigh_op_bnr_7')
// (13, 20, 'sp4_r_v_b_19')
// (13, 20, 'sp4_r_v_b_3')
// (13, 20, 'sp4_v_b_38')
// (13, 21, 'sp4_r_v_b_6')
// (13, 21, 'sp4_v_b_27')
// (13, 22, 'sp4_v_b_14')
// (13, 23, 'local_g1_3')
// (13, 23, 'lutff_7/in_1')
// (13, 23, 'sp4_v_b_3')
// (14, 16, 'sp4_v_t_38')
// (14, 17, 'local_g2_6')
// (14, 17, 'lutff_2/in_2')
// (14, 17, 'sp4_v_b_38')
// (14, 17, 'sp4_v_t_43')
// (14, 18, 'neigh_op_top_7')
// (14, 18, 'sp4_v_b_27')
// (14, 18, 'sp4_v_b_43')
// (14, 19, 'local_g1_7')
// (14, 19, 'lutff_7/in_1')
// (14, 19, 'lutff_7/out')
// (14, 19, 'sp12_h_r_6')
// (14, 19, 'sp4_h_r_14')
// (14, 19, 'sp4_v_b_14')
// (14, 19, 'sp4_v_b_30')
// (14, 20, 'neigh_op_bot_7')
// (14, 20, 'sp4_v_b_19')
// (14, 20, 'sp4_v_b_3')
// (14, 21, 'sp4_h_r_0')
// (14, 21, 'sp4_v_b_6')
// (15, 18, 'neigh_op_tnl_7')
// (15, 19, 'neigh_op_lft_7')
// (15, 19, 'sp12_h_r_9')
// (15, 19, 'sp4_h_r_27')
// (15, 20, 'neigh_op_bnl_7')
// (15, 21, 'local_g0_5')
// (15, 21, 'lutff_7/in_2')
// (15, 21, 'sp4_h_r_13')
// (16, 19, 'sp12_h_r_10')
// (16, 19, 'sp4_h_r_38')
// (16, 21, 'sp4_h_r_24')
// (17, 19, 'sp12_h_r_13')
// (17, 19, 'sp4_h_l_38')
// (17, 21, 'sp4_h_r_37')
// (17, 22, 'sp4_r_v_b_40')
// (17, 23, 'local_g1_5')
// (17, 23, 'lutff_7/in_1')
// (17, 23, 'sp4_r_v_b_29')
// (17, 24, 'sp4_r_v_b_16')
// (17, 25, 'sp4_r_v_b_5')
// (18, 19, 'sp12_h_r_14')
// (18, 21, 'sp4_h_l_37')
// (18, 21, 'sp4_v_t_40')
// (18, 22, 'sp4_v_b_40')
// (18, 23, 'sp4_v_b_29')
// (18, 24, 'sp4_v_b_16')
// (18, 25, 'sp4_v_b_5')
// (19, 19, 'sp12_h_r_17')
// (20, 19, 'sp12_h_r_18')
// (21, 19, 'sp12_h_r_21')
// (22, 19, 'sp12_h_r_22')
// (23, 19, 'sp12_h_l_22')

reg n514 = 0;
// (11, 19, 'local_g0_3')
// (11, 19, 'lutff_3/in_2')
// (11, 19, 'sp4_h_r_3')
// (11, 22, 'sp4_h_r_7')
// (12, 19, 'sp4_h_r_14')
// (12, 20, 'sp4_r_v_b_40')
// (12, 21, 'sp4_r_v_b_29')
// (12, 22, 'local_g0_2')
// (12, 22, 'lutff_3/in_1')
// (12, 22, 'sp4_h_r_18')
// (12, 22, 'sp4_r_v_b_16')
// (12, 23, 'sp4_r_v_b_5')
// (13, 16, 'sp4_r_v_b_43')
// (13, 17, 'local_g0_6')
// (13, 17, 'lutff_2/in_2')
// (13, 17, 'sp4_r_v_b_30')
// (13, 18, 'neigh_op_tnr_3')
// (13, 18, 'sp4_r_v_b_19')
// (13, 19, 'local_g3_3')
// (13, 19, 'lutff_3/in_3')
// (13, 19, 'neigh_op_rgt_3')
// (13, 19, 'sp4_h_r_11')
// (13, 19, 'sp4_h_r_27')
// (13, 19, 'sp4_r_v_b_6')
// (13, 19, 'sp4_v_t_40')
// (13, 20, 'neigh_op_bnr_3')
// (13, 20, 'sp4_v_b_40')
// (13, 21, 'sp4_v_b_29')
// (13, 22, 'sp4_h_r_31')
// (13, 22, 'sp4_v_b_16')
// (13, 23, 'local_g1_5')
// (13, 23, 'lutff_3/in_1')
// (13, 23, 'sp4_v_b_5')
// (14, 15, 'sp4_v_t_43')
// (14, 16, 'sp4_v_b_43')
// (14, 17, 'sp4_v_b_30')
// (14, 18, 'neigh_op_top_3')
// (14, 18, 'sp4_v_b_19')
// (14, 19, 'local_g1_3')
// (14, 19, 'lutff_3/in_1')
// (14, 19, 'lutff_3/out')
// (14, 19, 'sp4_h_r_22')
// (14, 19, 'sp4_h_r_38')
// (14, 19, 'sp4_r_v_b_39')
// (14, 19, 'sp4_v_b_6')
// (14, 20, 'neigh_op_bot_3')
// (14, 20, 'sp4_r_v_b_26')
// (14, 21, 'sp4_r_v_b_15')
// (14, 22, 'sp4_h_r_42')
// (14, 22, 'sp4_r_v_b_2')
// (15, 18, 'neigh_op_tnl_3')
// (15, 18, 'sp4_v_t_39')
// (15, 19, 'neigh_op_lft_3')
// (15, 19, 'sp4_h_l_38')
// (15, 19, 'sp4_h_r_35')
// (15, 19, 'sp4_v_b_39')
// (15, 20, 'neigh_op_bnl_3')
// (15, 20, 'sp4_v_b_26')
// (15, 21, 'local_g0_7')
// (15, 21, 'lutff_3/in_2')
// (15, 21, 'sp4_v_b_15')
// (15, 22, 'sp4_h_l_42')
// (15, 22, 'sp4_v_b_2')
// (16, 19, 'sp4_h_r_46')
// (16, 20, 'sp4_r_v_b_41')
// (16, 21, 'sp4_r_v_b_28')
// (16, 22, 'sp4_r_v_b_17')
// (16, 23, 'sp4_r_v_b_4')
// (17, 19, 'sp4_h_l_46')
// (17, 19, 'sp4_v_t_41')
// (17, 20, 'sp4_v_b_41')
// (17, 21, 'sp4_v_b_28')
// (17, 22, 'sp4_v_b_17')
// (17, 23, 'local_g1_4')
// (17, 23, 'lutff_3/in_2')
// (17, 23, 'sp4_v_b_4')

reg n515 = 0;
// (11, 19, 'local_g0_7')
// (11, 19, 'lutff_5/in_2')
// (11, 19, 'sp4_h_r_7')
// (12, 19, 'sp4_h_r_18')
// (12, 20, 'sp4_r_v_b_43')
// (12, 21, 'sp4_r_v_b_30')
// (12, 22, 'local_g3_3')
// (12, 22, 'lutff_5/in_1')
// (12, 22, 'sp4_r_v_b_19')
// (12, 23, 'sp4_r_v_b_6')
// (13, 16, 'sp4_r_v_b_47')
// (13, 17, 'sp4_r_v_b_34')
// (13, 18, 'neigh_op_tnr_5')
// (13, 18, 'sp4_r_v_b_23')
// (13, 19, 'local_g3_5')
// (13, 19, 'lutff_5/in_3')
// (13, 19, 'neigh_op_rgt_5')
// (13, 19, 'sp12_h_r_1')
// (13, 19, 'sp4_h_r_0')
// (13, 19, 'sp4_h_r_31')
// (13, 19, 'sp4_r_v_b_10')
// (13, 19, 'sp4_v_t_43')
// (13, 20, 'neigh_op_bnr_5')
// (13, 20, 'sp4_v_b_43')
// (13, 21, 'sp4_v_b_30')
// (13, 22, 'sp4_v_b_19')
// (13, 23, 'local_g0_6')
// (13, 23, 'lutff_5/in_1')
// (13, 23, 'sp4_v_b_6')
// (14, 15, 'sp4_v_t_47')
// (14, 16, 'sp4_v_b_47')
// (14, 17, 'local_g3_2')
// (14, 17, 'lutff_2/in_1')
// (14, 17, 'sp4_v_b_34')
// (14, 18, 'neigh_op_top_5')
// (14, 18, 'sp4_v_b_23')
// (14, 19, 'local_g1_5')
// (14, 19, 'lutff_5/in_1')
// (14, 19, 'lutff_5/out')
// (14, 19, 'sp12_h_r_2')
// (14, 19, 'sp4_h_r_13')
// (14, 19, 'sp4_h_r_42')
// (14, 19, 'sp4_v_b_10')
// (14, 20, 'neigh_op_bot_5')
// (14, 20, 'sp4_r_v_b_42')
// (14, 21, 'sp4_r_v_b_31')
// (14, 22, 'sp4_r_v_b_18')
// (14, 23, 'sp4_r_v_b_7')
// (15, 18, 'neigh_op_tnl_5')
// (15, 19, 'neigh_op_lft_5')
// (15, 19, 'sp12_h_r_5')
// (15, 19, 'sp4_h_l_42')
// (15, 19, 'sp4_h_r_24')
// (15, 19, 'sp4_v_t_42')
// (15, 20, 'neigh_op_bnl_5')
// (15, 20, 'sp4_v_b_42')
// (15, 21, 'local_g2_7')
// (15, 21, 'lutff_5/in_2')
// (15, 21, 'sp4_v_b_31')
// (15, 22, 'sp4_v_b_18')
// (15, 23, 'sp4_h_r_7')
// (15, 23, 'sp4_v_b_7')
// (16, 19, 'sp12_h_r_6')
// (16, 19, 'sp4_h_r_37')
// (16, 23, 'sp4_h_r_18')
// (17, 19, 'sp12_h_r_9')
// (17, 19, 'sp4_h_l_37')
// (17, 23, 'local_g3_7')
// (17, 23, 'lutff_5/in_1')
// (17, 23, 'sp4_h_r_31')
// (18, 19, 'sp12_h_r_10')
// (18, 23, 'sp4_h_r_42')
// (19, 19, 'sp12_h_r_13')
// (19, 23, 'sp4_h_l_42')
// (20, 19, 'sp12_h_r_14')
// (21, 19, 'sp12_h_r_17')
// (22, 19, 'sp12_h_r_18')
// (23, 19, 'sp12_h_r_21')
// (24, 19, 'sp12_h_r_22')
// (25, 19, 'sp12_h_l_22')

reg n516 = 0;
// (11, 19, 'local_g1_1')
// (11, 19, 'lutff_2/in_2')
// (11, 19, 'sp4_h_r_1')
// (11, 22, 'sp4_h_r_5')
// (12, 19, 'sp4_h_r_12')
// (12, 22, 'local_g0_0')
// (12, 22, 'lutff_2/in_2')
// (12, 22, 'sp4_h_r_16')
// (13, 16, 'sp4_r_v_b_41')
// (13, 17, 'local_g0_4')
// (13, 17, 'lutff_2/in_0')
// (13, 17, 'sp4_r_v_b_28')
// (13, 18, 'neigh_op_tnr_2')
// (13, 18, 'sp4_r_v_b_17')
// (13, 19, 'local_g3_2')
// (13, 19, 'lutff_2/in_3')
// (13, 19, 'neigh_op_rgt_2')
// (13, 19, 'sp4_h_r_25')
// (13, 19, 'sp4_h_r_9')
// (13, 19, 'sp4_r_v_b_4')
// (13, 20, 'neigh_op_bnr_2')
// (13, 20, 'sp4_r_v_b_42')
// (13, 21, 'sp4_r_v_b_31')
// (13, 22, 'sp4_h_r_29')
// (13, 22, 'sp4_r_v_b_18')
// (13, 23, 'local_g1_7')
// (13, 23, 'lutff_2/in_2')
// (13, 23, 'sp4_r_v_b_7')
// (14, 15, 'sp4_v_t_41')
// (14, 16, 'sp4_v_b_41')
// (14, 17, 'sp4_v_b_28')
// (14, 18, 'neigh_op_top_2')
// (14, 18, 'sp4_v_b_17')
// (14, 19, 'local_g1_4')
// (14, 19, 'lutff_2/in_1')
// (14, 19, 'lutff_2/out')
// (14, 19, 'sp4_h_r_20')
// (14, 19, 'sp4_h_r_36')
// (14, 19, 'sp4_r_v_b_37')
// (14, 19, 'sp4_v_b_4')
// (14, 19, 'sp4_v_t_42')
// (14, 20, 'neigh_op_bot_2')
// (14, 20, 'sp4_r_v_b_24')
// (14, 20, 'sp4_v_b_42')
// (14, 21, 'sp4_r_v_b_13')
// (14, 21, 'sp4_v_b_31')
// (14, 22, 'sp4_h_r_40')
// (14, 22, 'sp4_r_v_b_0')
// (14, 22, 'sp4_v_b_18')
// (14, 23, 'sp4_v_b_7')
// (15, 18, 'neigh_op_tnl_2')
// (15, 18, 'sp4_v_t_37')
// (15, 19, 'neigh_op_lft_2')
// (15, 19, 'sp4_h_l_36')
// (15, 19, 'sp4_h_r_33')
// (15, 19, 'sp4_v_b_37')
// (15, 20, 'neigh_op_bnl_2')
// (15, 20, 'sp4_v_b_24')
// (15, 21, 'local_g1_5')
// (15, 21, 'lutff_2/in_2')
// (15, 21, 'sp4_v_b_13')
// (15, 22, 'sp4_h_l_40')
// (15, 22, 'sp4_v_b_0')
// (16, 19, 'sp4_h_r_44')
// (16, 20, 'sp4_r_v_b_44')
// (16, 21, 'sp4_r_v_b_33')
// (16, 22, 'sp4_r_v_b_20')
// (16, 23, 'sp4_r_v_b_9')
// (17, 19, 'sp4_h_l_44')
// (17, 19, 'sp4_v_t_44')
// (17, 20, 'sp4_v_b_44')
// (17, 21, 'sp4_v_b_33')
// (17, 22, 'sp4_v_b_20')
// (17, 23, 'local_g0_1')
// (17, 23, 'lutff_2/in_1')
// (17, 23, 'sp4_v_b_9')

wire n517;
// (11, 19, 'lutff_7/cout')
// (11, 20, 'carry_in')
// (11, 20, 'carry_in_mux')

reg n518 = 0;
// (11, 19, 'neigh_op_tnr_0')
// (11, 20, 'neigh_op_rgt_0')
// (11, 21, 'neigh_op_bnr_0')
// (12, 19, 'neigh_op_top_0')
// (12, 20, 'lutff_0/out')
// (12, 21, 'local_g0_0')
// (12, 21, 'lutff_0/in_0')
// (12, 21, 'neigh_op_bot_0')
// (13, 19, 'neigh_op_tnl_0')
// (13, 20, 'neigh_op_lft_0')
// (13, 21, 'neigh_op_bnl_0')

reg n519 = 0;
// (11, 19, 'neigh_op_tnr_2')
// (11, 20, 'neigh_op_rgt_2')
// (11, 21, 'neigh_op_bnr_2')
// (12, 19, 'neigh_op_top_2')
// (12, 20, 'lutff_2/out')
// (12, 21, 'local_g1_2')
// (12, 21, 'lutff_2/in_3')
// (12, 21, 'neigh_op_bot_2')
// (13, 19, 'neigh_op_tnl_2')
// (13, 20, 'neigh_op_lft_2')
// (13, 21, 'neigh_op_bnl_2')

reg n520 = 0;
// (11, 19, 'neigh_op_tnr_3')
// (11, 20, 'neigh_op_rgt_3')
// (11, 21, 'neigh_op_bnr_3')
// (12, 19, 'neigh_op_top_3')
// (12, 20, 'lutff_3/out')
// (12, 21, 'local_g0_3')
// (12, 21, 'lutff_3/in_0')
// (12, 21, 'neigh_op_bot_3')
// (13, 19, 'neigh_op_tnl_3')
// (13, 20, 'neigh_op_lft_3')
// (13, 21, 'neigh_op_bnl_3')

reg n521 = 0;
// (11, 19, 'neigh_op_tnr_5')
// (11, 20, 'neigh_op_rgt_5')
// (11, 21, 'neigh_op_bnr_5')
// (12, 19, 'neigh_op_top_5')
// (12, 20, 'lutff_5/out')
// (12, 21, 'local_g0_5')
// (12, 21, 'lutff_5/in_0')
// (12, 21, 'neigh_op_bot_5')
// (13, 19, 'neigh_op_tnl_5')
// (13, 20, 'neigh_op_lft_5')
// (13, 21, 'neigh_op_bnl_5')

reg n522 = 0;
// (11, 19, 'neigh_op_tnr_6')
// (11, 20, 'neigh_op_rgt_6')
// (11, 21, 'neigh_op_bnr_6')
// (12, 19, 'neigh_op_top_6')
// (12, 20, 'lutff_6/out')
// (12, 21, 'local_g0_6')
// (12, 21, 'lutff_6/in_0')
// (12, 21, 'neigh_op_bot_6')
// (13, 19, 'neigh_op_tnl_6')
// (13, 20, 'neigh_op_lft_6')
// (13, 21, 'neigh_op_bnl_6')

reg n523 = 0;
// (11, 19, 'neigh_op_tnr_7')
// (11, 20, 'neigh_op_rgt_7')
// (11, 21, 'neigh_op_bnr_7')
// (12, 19, 'neigh_op_top_7')
// (12, 20, 'lutff_7/out')
// (12, 21, 'local_g1_7')
// (12, 21, 'lutff_7/in_3')
// (12, 21, 'neigh_op_bot_7')
// (13, 19, 'neigh_op_tnl_7')
// (13, 20, 'neigh_op_lft_7')
// (13, 21, 'neigh_op_bnl_7')

wire n524;
// (11, 19, 'sp12_h_r_0')
// (12, 18, 'neigh_op_tnr_6')
// (12, 19, 'neigh_op_rgt_6')
// (12, 19, 'sp12_h_r_3')
// (12, 20, 'neigh_op_bnr_6')
// (13, 18, 'neigh_op_top_6')
// (13, 19, 'local_g2_6')
// (13, 19, 'lutff_6/in_2')
// (13, 19, 'lutff_6/out')
// (13, 19, 'sp12_h_r_4')
// (13, 20, 'neigh_op_bot_6')
// (14, 18, 'neigh_op_tnl_6')
// (14, 19, 'neigh_op_lft_6')
// (14, 19, 'sp12_h_r_7')
// (14, 20, 'neigh_op_bnl_6')
// (15, 19, 'sp12_h_r_8')
// (16, 19, 'sp12_h_r_11')
// (17, 19, 'local_g0_4')
// (17, 19, 'lutff_6/in_2')
// (17, 19, 'sp12_h_r_12')
// (18, 19, 'sp12_h_r_15')
// (19, 19, 'sp12_h_r_16')
// (20, 19, 'sp12_h_r_19')
// (21, 19, 'sp12_h_r_20')
// (22, 19, 'sp12_h_r_23')
// (23, 19, 'sp12_h_l_23')

wire n525;
// (11, 19, 'sp4_r_v_b_44')
// (11, 20, 'sp4_r_v_b_33')
// (11, 21, 'local_g3_4')
// (11, 21, 'lutff_3/in_0')
// (11, 21, 'sp4_r_v_b_20')
// (11, 22, 'sp4_r_v_b_9')
// (12, 12, 'sp12_h_r_0')
// (12, 18, 'sp4_h_r_9')
// (12, 18, 'sp4_v_t_44')
// (12, 19, 'sp4_v_b_44')
// (12, 20, 'sp4_v_b_33')
// (12, 21, 'sp4_v_b_20')
// (12, 22, 'sp4_v_b_9')
// (13, 12, 'sp12_h_r_3')
// (13, 18, 'sp4_h_r_20')
// (14, 12, 'sp12_h_r_4')
// (14, 18, 'sp4_h_r_33')
// (15, 11, 'neigh_op_tnr_0')
// (15, 11, 'sp4_r_v_b_45')
// (15, 12, 'neigh_op_rgt_0')
// (15, 12, 'sp12_h_r_7')
// (15, 12, 'sp4_r_v_b_32')
// (15, 13, 'neigh_op_bnr_0')
// (15, 13, 'sp4_r_v_b_21')
// (15, 14, 'local_g2_0')
// (15, 14, 'lutff_1/in_1')
// (15, 14, 'sp4_r_v_b_8')
// (15, 15, 'sp4_r_v_b_41')
// (15, 16, 'local_g0_4')
// (15, 16, 'local_g1_4')
// (15, 16, 'lutff_1/in_0')
// (15, 16, 'lutff_2/in_0')
// (15, 16, 'sp4_r_v_b_28')
// (15, 17, 'sp4_r_v_b_17')
// (15, 18, 'sp4_h_r_44')
// (15, 18, 'sp4_r_v_b_4')
// (16, 8, 'sp12_v_t_23')
// (16, 9, 'sp12_v_b_23')
// (16, 10, 'sp12_v_b_20')
// (16, 10, 'sp4_v_t_45')
// (16, 11, 'neigh_op_top_0')
// (16, 11, 'sp12_v_b_19')
// (16, 11, 'sp4_v_b_45')
// (16, 12, 'local_g0_0')
// (16, 12, 'lutff_0/out')
// (16, 12, 'lutff_3/in_1')
// (16, 12, 'sp12_h_r_8')
// (16, 12, 'sp12_v_b_16')
// (16, 12, 'sp4_v_b_32')
// (16, 13, 'neigh_op_bot_0')
// (16, 13, 'sp12_v_b_15')
// (16, 13, 'sp4_v_b_21')
// (16, 14, 'local_g0_0')
// (16, 14, 'lutff_2/in_0')
// (16, 14, 'lutff_6/in_0')
// (16, 14, 'lutff_7/in_1')
// (16, 14, 'sp12_v_b_12')
// (16, 14, 'sp4_v_b_8')
// (16, 14, 'sp4_v_t_41')
// (16, 15, 'local_g3_3')
// (16, 15, 'lutff_5/in_1')
// (16, 15, 'sp12_v_b_11')
// (16, 15, 'sp4_v_b_41')
// (16, 16, 'sp12_v_b_8')
// (16, 16, 'sp4_v_b_28')
// (16, 17, 'sp12_v_b_7')
// (16, 17, 'sp4_v_b_17')
// (16, 18, 'sp12_v_b_4')
// (16, 18, 'sp4_h_l_44')
// (16, 18, 'sp4_v_b_4')
// (16, 19, 'sp12_v_b_3')
// (16, 20, 'local_g2_0')
// (16, 20, 'lutff_7/in_1')
// (16, 20, 'sp12_v_b_0')
// (17, 11, 'neigh_op_tnl_0')
// (17, 12, 'neigh_op_lft_0')
// (17, 12, 'sp12_h_r_11')
// (17, 13, 'neigh_op_bnl_0')
// (18, 12, 'sp12_h_r_12')
// (19, 12, 'local_g1_7')
// (19, 12, 'lutff_1/in_1')
// (19, 12, 'sp12_h_r_15')
// (19, 12, 'sp4_h_r_9')
// (20, 12, 'sp12_h_r_16')
// (20, 12, 'sp4_h_r_20')
// (21, 12, 'sp12_h_r_19')
// (21, 12, 'sp4_h_r_33')
// (22, 12, 'sp12_h_r_20')
// (22, 12, 'sp4_h_r_44')
// (22, 13, 'sp4_r_v_b_44')
// (22, 14, 'sp4_r_v_b_33')
// (22, 15, 'local_g3_4')
// (22, 15, 'lutff_0/in_1')
// (22, 15, 'lutff_5/in_2')
// (22, 15, 'lutff_6/in_1')
// (22, 15, 'lutff_7/in_2')
// (22, 15, 'sp4_r_v_b_20')
// (22, 16, 'sp4_r_v_b_9')
// (23, 12, 'sp12_h_r_23')
// (23, 12, 'sp4_h_l_44')
// (23, 12, 'sp4_v_t_44')
// (23, 13, 'sp4_v_b_44')
// (23, 14, 'sp4_v_b_33')
// (23, 15, 'sp4_v_b_20')
// (23, 16, 'sp4_v_b_9')
// (24, 12, 'sp12_h_l_23')

reg n526 = 0;
// (11, 20, 'local_g0_1')
// (11, 20, 'lutff_7/in_2')
// (11, 20, 'sp12_h_r_1')
// (12, 20, 'sp12_h_r_2')
// (12, 21, 'sp4_r_v_b_38')
// (12, 22, 'sp4_r_v_b_27')
// (12, 23, 'local_g2_6')
// (12, 23, 'lutff_7/in_1')
// (12, 23, 'sp4_r_v_b_14')
// (12, 24, 'sp4_r_v_b_3')
// (13, 18, 'sp4_r_v_b_38')
// (13, 19, 'neigh_op_tnr_7')
// (13, 19, 'sp4_r_v_b_27')
// (13, 20, 'local_g2_7')
// (13, 20, 'lutff_7/in_0')
// (13, 20, 'neigh_op_rgt_7')
// (13, 20, 'sp12_h_r_5')
// (13, 20, 'sp4_h_r_3')
// (13, 20, 'sp4_r_v_b_14')
// (13, 20, 'sp4_v_t_38')
// (13, 21, 'neigh_op_bnr_7')
// (13, 21, 'sp4_r_v_b_3')
// (13, 21, 'sp4_v_b_38')
// (13, 22, 'sp4_r_v_b_43')
// (13, 22, 'sp4_v_b_27')
// (13, 23, 'sp4_r_v_b_30')
// (13, 23, 'sp4_v_b_14')
// (13, 24, 'local_g3_3')
// (13, 24, 'lutff_7/in_1')
// (13, 24, 'sp4_r_v_b_19')
// (13, 24, 'sp4_v_b_3')
// (13, 25, 'sp4_r_v_b_6')
// (14, 17, 'local_g0_0')
// (14, 17, 'lutff_0/in_2')
// (14, 17, 'sp4_h_r_8')
// (14, 17, 'sp4_v_t_38')
// (14, 18, 'sp4_v_b_38')
// (14, 19, 'neigh_op_top_7')
// (14, 19, 'sp4_v_b_27')
// (14, 20, 'local_g1_7')
// (14, 20, 'lutff_7/in_1')
// (14, 20, 'lutff_7/out')
// (14, 20, 'sp12_h_r_6')
// (14, 20, 'sp4_h_r_14')
// (14, 20, 'sp4_r_v_b_47')
// (14, 20, 'sp4_v_b_14')
// (14, 21, 'neigh_op_bot_7')
// (14, 21, 'sp4_r_v_b_34')
// (14, 21, 'sp4_v_b_3')
// (14, 21, 'sp4_v_t_43')
// (14, 22, 'sp4_r_v_b_23')
// (14, 22, 'sp4_v_b_43')
// (14, 23, 'sp4_r_v_b_10')
// (14, 23, 'sp4_v_b_30')
// (14, 24, 'sp4_v_b_19')
// (14, 25, 'sp4_v_b_6')
// (15, 17, 'sp4_h_r_21')
// (15, 19, 'neigh_op_tnl_7')
// (15, 19, 'sp4_v_t_47')
// (15, 20, 'neigh_op_lft_7')
// (15, 20, 'sp12_h_r_9')
// (15, 20, 'sp4_h_r_27')
// (15, 20, 'sp4_v_b_47')
// (15, 21, 'neigh_op_bnl_7')
// (15, 21, 'sp4_v_b_34')
// (15, 22, 'local_g0_7')
// (15, 22, 'lutff_7/in_2')
// (15, 22, 'sp4_v_b_23')
// (15, 23, 'sp4_v_b_10')
// (16, 17, 'sp4_h_r_32')
// (16, 20, 'sp12_h_r_10')
// (16, 20, 'sp4_h_r_38')
// (16, 21, 'sp4_r_v_b_45')
// (16, 22, 'sp4_r_v_b_32')
// (16, 23, 'sp4_r_v_b_21')
// (16, 24, 'sp4_r_v_b_8')
// (17, 17, 'sp4_h_r_45')
// (17, 20, 'local_g0_5')
// (17, 20, 'lutff_7/in_0')
// (17, 20, 'sp12_h_r_13')
// (17, 20, 'sp4_h_l_38')
// (17, 20, 'sp4_v_t_45')
// (17, 21, 'sp4_v_b_45')
// (17, 22, 'sp4_v_b_32')
// (17, 23, 'sp4_v_b_21')
// (17, 24, 'local_g0_0')
// (17, 24, 'lutff_7/in_1')
// (17, 24, 'sp4_v_b_8')
// (18, 17, 'sp4_h_l_45')
// (18, 20, 'sp12_h_r_14')
// (19, 20, 'sp12_h_r_17')
// (20, 20, 'sp12_h_r_18')
// (21, 20, 'sp12_h_r_21')
// (22, 20, 'sp12_h_r_22')
// (23, 20, 'sp12_h_l_22')

reg n527 = 0;
// (11, 20, 'local_g0_3')
// (11, 20, 'lutff_3/in_2')
// (11, 20, 'sp4_h_r_3')
// (11, 23, 'sp4_h_r_2')
// (12, 20, 'sp4_h_r_14')
// (12, 21, 'sp4_r_v_b_46')
// (12, 22, 'sp4_r_v_b_35')
// (12, 23, 'local_g1_7')
// (12, 23, 'lutff_3/in_1')
// (12, 23, 'sp4_h_r_15')
// (12, 23, 'sp4_r_v_b_22')
// (12, 24, 'sp4_r_v_b_11')
// (13, 17, 'sp4_r_v_b_43')
// (13, 18, 'sp4_r_v_b_30')
// (13, 19, 'neigh_op_tnr_3')
// (13, 19, 'sp4_r_v_b_19')
// (13, 20, 'local_g3_3')
// (13, 20, 'lutff_3/in_3')
// (13, 20, 'neigh_op_rgt_3')
// (13, 20, 'sp4_h_r_11')
// (13, 20, 'sp4_h_r_27')
// (13, 20, 'sp4_r_v_b_6')
// (13, 20, 'sp4_v_t_46')
// (13, 21, 'neigh_op_bnr_3')
// (13, 21, 'sp4_v_b_46')
// (13, 22, 'sp4_v_b_35')
// (13, 23, 'sp4_h_r_26')
// (13, 23, 'sp4_v_b_22')
// (13, 24, 'local_g1_3')
// (13, 24, 'lutff_3/in_1')
// (13, 24, 'sp4_v_b_11')
// (14, 16, 'sp4_v_t_43')
// (14, 17, 'local_g3_3')
// (14, 17, 'lutff_0/in_0')
// (14, 17, 'sp4_v_b_43')
// (14, 18, 'sp4_v_b_30')
// (14, 19, 'neigh_op_top_3')
// (14, 19, 'sp4_v_b_19')
// (14, 20, 'local_g1_3')
// (14, 20, 'lutff_3/in_1')
// (14, 20, 'lutff_3/out')
// (14, 20, 'sp4_h_r_22')
// (14, 20, 'sp4_h_r_38')
// (14, 20, 'sp4_h_r_6')
// (14, 20, 'sp4_r_v_b_39')
// (14, 20, 'sp4_v_b_6')
// (14, 21, 'neigh_op_bot_3')
// (14, 21, 'sp4_r_v_b_26')
// (14, 22, 'sp4_r_v_b_15')
// (14, 23, 'sp4_h_r_39')
// (14, 23, 'sp4_r_v_b_2')
// (15, 19, 'neigh_op_tnl_3')
// (15, 19, 'sp4_v_t_39')
// (15, 20, 'neigh_op_lft_3')
// (15, 20, 'sp4_h_l_38')
// (15, 20, 'sp4_h_r_19')
// (15, 20, 'sp4_h_r_35')
// (15, 20, 'sp4_v_b_39')
// (15, 21, 'neigh_op_bnl_3')
// (15, 21, 'sp4_v_b_26')
// (15, 22, 'local_g1_7')
// (15, 22, 'lutff_3/in_1')
// (15, 22, 'sp4_v_b_15')
// (15, 23, 'sp4_h_l_39')
// (15, 23, 'sp4_v_b_2')
// (16, 20, 'sp4_h_r_30')
// (16, 20, 'sp4_h_r_46')
// (17, 20, 'local_g3_3')
// (17, 20, 'lutff_3/in_3')
// (17, 20, 'sp4_h_l_46')
// (17, 20, 'sp4_h_r_43')
// (17, 21, 'sp4_r_v_b_43')
// (17, 22, 'sp4_r_v_b_30')
// (17, 23, 'sp4_r_v_b_19')
// (17, 24, 'local_g1_6')
// (17, 24, 'lutff_3/in_2')
// (17, 24, 'sp4_r_v_b_6')
// (18, 20, 'sp4_h_l_43')
// (18, 20, 'sp4_v_t_43')
// (18, 21, 'sp4_v_b_43')
// (18, 22, 'sp4_v_b_30')
// (18, 23, 'sp4_v_b_19')
// (18, 24, 'sp4_v_b_6')

reg n528 = 0;
// (11, 20, 'local_g1_1')
// (11, 20, 'lutff_2/in_2')
// (11, 20, 'sp4_h_r_1')
// (11, 23, 'sp4_h_r_5')
// (12, 20, 'sp4_h_r_12')
// (12, 23, 'local_g0_0')
// (12, 23, 'lutff_2/in_2')
// (12, 23, 'sp4_h_r_16')
// (13, 17, 'sp4_r_v_b_41')
// (13, 18, 'sp4_r_v_b_28')
// (13, 19, 'neigh_op_tnr_2')
// (13, 19, 'sp4_r_v_b_17')
// (13, 20, 'local_g2_2')
// (13, 20, 'lutff_2/in_0')
// (13, 20, 'neigh_op_rgt_2')
// (13, 20, 'sp4_h_r_25')
// (13, 20, 'sp4_r_v_b_36')
// (13, 20, 'sp4_r_v_b_4')
// (13, 21, 'neigh_op_bnr_2')
// (13, 21, 'sp4_r_v_b_25')
// (13, 22, 'sp4_r_v_b_12')
// (13, 23, 'sp4_h_r_29')
// (13, 23, 'sp4_r_v_b_1')
// (13, 24, 'local_g3_1')
// (13, 24, 'lutff_2/in_2')
// (13, 24, 'sp4_r_v_b_41')
// (13, 25, 'sp4_r_v_b_28')
// (13, 26, 'sp4_r_v_b_17')
// (13, 27, 'sp4_r_v_b_4')
// (14, 16, 'sp4_v_t_41')
// (14, 17, 'local_g2_1')
// (14, 17, 'lutff_0/in_1')
// (14, 17, 'sp4_v_b_41')
// (14, 18, 'sp4_v_b_28')
// (14, 19, 'neigh_op_top_2')
// (14, 19, 'sp4_v_b_17')
// (14, 19, 'sp4_v_t_36')
// (14, 20, 'local_g1_2')
// (14, 20, 'lutff_2/in_1')
// (14, 20, 'lutff_2/out')
// (14, 20, 'sp4_h_r_36')
// (14, 20, 'sp4_h_r_4')
// (14, 20, 'sp4_r_v_b_37')
// (14, 20, 'sp4_v_b_36')
// (14, 20, 'sp4_v_b_4')
// (14, 21, 'neigh_op_bot_2')
// (14, 21, 'sp4_r_v_b_24')
// (14, 21, 'sp4_v_b_25')
// (14, 22, 'sp4_r_v_b_13')
// (14, 22, 'sp4_v_b_12')
// (14, 23, 'sp4_h_r_40')
// (14, 23, 'sp4_r_v_b_0')
// (14, 23, 'sp4_v_b_1')
// (14, 23, 'sp4_v_t_41')
// (14, 24, 'sp4_v_b_41')
// (14, 25, 'sp4_v_b_28')
// (14, 26, 'sp4_v_b_17')
// (14, 27, 'sp4_v_b_4')
// (15, 19, 'neigh_op_tnl_2')
// (15, 19, 'sp4_v_t_37')
// (15, 20, 'neigh_op_lft_2')
// (15, 20, 'sp4_h_l_36')
// (15, 20, 'sp4_h_r_17')
// (15, 20, 'sp4_v_b_37')
// (15, 21, 'neigh_op_bnl_2')
// (15, 21, 'sp4_v_b_24')
// (15, 22, 'local_g0_5')
// (15, 22, 'lutff_2/in_1')
// (15, 22, 'sp4_v_b_13')
// (15, 23, 'sp4_h_l_40')
// (15, 23, 'sp4_v_b_0')
// (16, 20, 'sp4_h_r_28')
// (17, 20, 'local_g2_1')
// (17, 20, 'lutff_2/in_3')
// (17, 20, 'sp4_h_r_41')
// (17, 21, 'sp4_r_v_b_41')
// (17, 22, 'sp4_r_v_b_28')
// (17, 23, 'sp4_r_v_b_17')
// (17, 24, 'local_g1_4')
// (17, 24, 'lutff_2/in_1')
// (17, 24, 'sp4_r_v_b_4')
// (18, 20, 'sp4_h_l_41')
// (18, 20, 'sp4_v_t_41')
// (18, 21, 'sp4_v_b_41')
// (18, 22, 'sp4_v_b_28')
// (18, 23, 'sp4_v_b_17')
// (18, 24, 'sp4_v_b_4')

wire n529;
// (11, 20, 'lutff_7/cout')
// (11, 21, 'carry_in')
// (11, 21, 'carry_in_mux')
// (11, 21, 'lutff_0/in_3')

wire n530;
// (11, 20, 'neigh_op_tnr_0')
// (11, 21, 'neigh_op_rgt_0')
// (11, 22, 'neigh_op_bnr_0')
// (12, 20, 'neigh_op_top_0')
// (12, 21, 'local_g3_0')
// (12, 21, 'lutff_0/in_1')
// (12, 21, 'lutff_0/out')
// (12, 22, 'neigh_op_bot_0')
// (13, 20, 'neigh_op_tnl_0')
// (13, 21, 'neigh_op_lft_0')
// (13, 22, 'neigh_op_bnl_0')

wire n531;
// (11, 20, 'neigh_op_tnr_1')
// (11, 21, 'neigh_op_rgt_1')
// (11, 22, 'neigh_op_bnr_1')
// (12, 20, 'neigh_op_top_1')
// (12, 21, 'local_g3_1')
// (12, 21, 'lutff_1/in_1')
// (12, 21, 'lutff_1/out')
// (12, 22, 'neigh_op_bot_1')
// (13, 20, 'neigh_op_tnl_1')
// (13, 21, 'neigh_op_lft_1')
// (13, 22, 'neigh_op_bnl_1')

wire n532;
// (11, 20, 'neigh_op_tnr_2')
// (11, 21, 'neigh_op_rgt_2')
// (11, 22, 'neigh_op_bnr_2')
// (12, 20, 'neigh_op_top_2')
// (12, 21, 'local_g2_2')
// (12, 21, 'lutff_2/in_2')
// (12, 21, 'lutff_2/out')
// (12, 22, 'neigh_op_bot_2')
// (13, 20, 'neigh_op_tnl_2')
// (13, 21, 'neigh_op_lft_2')
// (13, 22, 'neigh_op_bnl_2')

wire n533;
// (11, 20, 'neigh_op_tnr_3')
// (11, 21, 'neigh_op_rgt_3')
// (11, 22, 'neigh_op_bnr_3')
// (12, 20, 'neigh_op_top_3')
// (12, 21, 'local_g2_3')
// (12, 21, 'lutff_3/in_2')
// (12, 21, 'lutff_3/out')
// (12, 22, 'neigh_op_bot_3')
// (13, 20, 'neigh_op_tnl_3')
// (13, 21, 'neigh_op_lft_3')
// (13, 22, 'neigh_op_bnl_3')

wire n534;
// (11, 20, 'neigh_op_tnr_4')
// (11, 21, 'neigh_op_rgt_4')
// (11, 22, 'neigh_op_bnr_4')
// (12, 20, 'neigh_op_top_4')
// (12, 21, 'local_g3_4')
// (12, 21, 'lutff_4/in_1')
// (12, 21, 'lutff_4/out')
// (12, 22, 'neigh_op_bot_4')
// (13, 20, 'neigh_op_tnl_4')
// (13, 21, 'neigh_op_lft_4')
// (13, 22, 'neigh_op_bnl_4')

wire n535;
// (11, 20, 'neigh_op_tnr_5')
// (11, 21, 'neigh_op_rgt_5')
// (11, 22, 'neigh_op_bnr_5')
// (12, 20, 'neigh_op_top_5')
// (12, 21, 'local_g3_5')
// (12, 21, 'lutff_5/in_1')
// (12, 21, 'lutff_5/out')
// (12, 22, 'neigh_op_bot_5')
// (13, 20, 'neigh_op_tnl_5')
// (13, 21, 'neigh_op_lft_5')
// (13, 22, 'neigh_op_bnl_5')

wire n536;
// (11, 20, 'neigh_op_tnr_6')
// (11, 21, 'neigh_op_rgt_6')
// (11, 22, 'neigh_op_bnr_6')
// (12, 20, 'neigh_op_top_6')
// (12, 21, 'local_g1_6')
// (12, 21, 'lutff_6/in_1')
// (12, 21, 'lutff_6/out')
// (12, 22, 'neigh_op_bot_6')
// (13, 20, 'neigh_op_tnl_6')
// (13, 21, 'neigh_op_lft_6')
// (13, 22, 'neigh_op_bnl_6')

wire n537;
// (11, 20, 'neigh_op_tnr_7')
// (11, 21, 'neigh_op_rgt_7')
// (11, 22, 'neigh_op_bnr_7')
// (12, 20, 'neigh_op_top_7')
// (12, 21, 'local_g3_7')
// (12, 21, 'lutff_7/in_1')
// (12, 21, 'lutff_7/out')
// (12, 22, 'neigh_op_bot_7')
// (13, 20, 'neigh_op_tnl_7')
// (13, 21, 'neigh_op_lft_7')
// (13, 22, 'neigh_op_bnl_7')

wire n538;
// (11, 20, 'sp4_r_v_b_43')
// (11, 21, 'sp4_r_v_b_30')
// (11, 22, 'sp4_r_v_b_19')
// (11, 23, 'sp4_r_v_b_6')
// (12, 19, 'sp4_h_r_6')
// (12, 19, 'sp4_v_t_43')
// (12, 20, 'local_g3_3')
// (12, 20, 'lutff_global/cen')
// (12, 20, 'sp4_v_b_43')
// (12, 21, 'sp4_v_b_30')
// (12, 22, 'sp4_v_b_19')
// (12, 23, 'sp4_h_r_2')
// (12, 23, 'sp4_v_b_6')
// (13, 19, 'sp4_h_r_19')
// (13, 23, 'sp4_h_r_15')
// (14, 19, 'sp4_h_r_30')
// (14, 23, 'local_g2_2')
// (14, 23, 'lutff_global/cen')
// (14, 23, 'sp4_h_r_26')
// (15, 11, 'neigh_op_tnr_4')
// (15, 12, 'neigh_op_rgt_4')
// (15, 12, 'sp4_r_v_b_40')
// (15, 13, 'neigh_op_bnr_4')
// (15, 13, 'sp4_r_v_b_29')
// (15, 14, 'sp4_r_v_b_16')
// (15, 15, 'sp4_r_v_b_5')
// (15, 16, 'sp4_r_v_b_36')
// (15, 17, 'sp4_r_v_b_25')
// (15, 18, 'sp4_r_v_b_12')
// (15, 19, 'sp4_h_r_43')
// (15, 19, 'sp4_r_v_b_1')
// (15, 20, 'sp4_r_v_b_44')
// (15, 21, 'sp4_r_v_b_33')
// (15, 22, 'sp4_r_v_b_20')
// (15, 23, 'sp4_h_r_39')
// (15, 23, 'sp4_r_v_b_9')
// (16, 11, 'neigh_op_top_4')
// (16, 11, 'sp4_v_t_40')
// (16, 12, 'lutff_4/out')
// (16, 12, 'sp4_v_b_40')
// (16, 13, 'neigh_op_bot_4')
// (16, 13, 'sp4_v_b_29')
// (16, 14, 'sp4_v_b_16')
// (16, 15, 'sp4_v_b_5')
// (16, 15, 'sp4_v_t_36')
// (16, 16, 'sp4_v_b_36')
// (16, 17, 'sp4_v_b_25')
// (16, 18, 'sp4_v_b_12')
// (16, 19, 'sp4_h_l_43')
// (16, 19, 'sp4_v_b_1')
// (16, 19, 'sp4_v_t_44')
// (16, 20, 'sp4_v_b_44')
// (16, 21, 'sp4_v_b_33')
// (16, 22, 'sp4_v_b_20')
// (16, 23, 'sp4_h_l_39')
// (16, 23, 'sp4_v_b_9')
// (17, 11, 'neigh_op_tnl_4')
// (17, 12, 'neigh_op_lft_4')
// (17, 13, 'neigh_op_bnl_4')

reg n539 = 0;
// (11, 20, 'sp4_r_v_b_46')
// (11, 21, 'sp4_r_v_b_35')
// (11, 22, 'sp4_r_v_b_22')
// (11, 23, 'sp4_r_v_b_11')
// (12, 19, 'sp4_v_t_46')
// (12, 20, 'sp4_v_b_46')
// (12, 21, 'local_g3_3')
// (12, 21, 'lutff_1/in_3')
// (12, 21, 'sp4_v_b_35')
// (12, 22, 'sp4_v_b_22')
// (12, 23, 'sp4_h_r_6')
// (12, 23, 'sp4_v_b_11')
// (13, 22, 'neigh_op_tnr_7')
// (13, 23, 'neigh_op_rgt_7')
// (13, 23, 'sp4_h_r_19')
// (13, 24, 'neigh_op_bnr_7')
// (14, 22, 'neigh_op_top_7')
// (14, 23, 'lutff_7/out')
// (14, 23, 'sp4_h_r_30')
// (14, 24, 'neigh_op_bot_7')
// (15, 22, 'neigh_op_tnl_7')
// (15, 23, 'neigh_op_lft_7')
// (15, 23, 'sp4_h_r_43')
// (15, 24, 'neigh_op_bnl_7')
// (16, 23, 'sp4_h_l_43')

wire n540;
// (11, 21, 'local_g1_3')
// (11, 21, 'lutff_3/in_3')
// (11, 21, 'sp4_h_r_3')
// (12, 21, 'sp4_h_r_14')
// (13, 21, 'sp4_h_r_27')
// (14, 13, 'neigh_op_tnr_3')
// (14, 14, 'neigh_op_rgt_3')
// (14, 14, 'sp4_r_v_b_38')
// (14, 15, 'neigh_op_bnr_3')
// (14, 15, 'sp4_r_v_b_27')
// (14, 16, 'sp4_r_v_b_14')
// (14, 17, 'sp4_r_v_b_3')
// (14, 18, 'sp4_r_v_b_38')
// (14, 19, 'sp4_r_v_b_27')
// (14, 20, 'sp4_r_v_b_14')
// (14, 21, 'sp4_h_r_38')
// (14, 21, 'sp4_r_v_b_3')
// (15, 13, 'neigh_op_top_3')
// (15, 13, 'sp4_v_t_38')
// (15, 14, 'local_g1_3')
// (15, 14, 'lutff_1/in_3')
// (15, 14, 'lutff_3/out')
// (15, 14, 'sp4_r_v_b_39')
// (15, 14, 'sp4_v_b_38')
// (15, 15, 'neigh_op_bot_3')
// (15, 15, 'sp4_r_v_b_26')
// (15, 15, 'sp4_v_b_27')
// (15, 16, 'local_g1_6')
// (15, 16, 'lutff_6/in_3')
// (15, 16, 'sp4_r_v_b_15')
// (15, 16, 'sp4_v_b_14')
// (15, 17, 'sp4_r_v_b_2')
// (15, 17, 'sp4_v_b_3')
// (15, 17, 'sp4_v_t_38')
// (15, 18, 'sp4_r_v_b_39')
// (15, 18, 'sp4_v_b_38')
// (15, 19, 'sp4_r_v_b_26')
// (15, 19, 'sp4_v_b_27')
// (15, 20, 'sp4_r_v_b_15')
// (15, 20, 'sp4_v_b_14')
// (15, 21, 'sp4_h_l_38')
// (15, 21, 'sp4_r_v_b_2')
// (15, 21, 'sp4_v_b_3')
// (16, 13, 'neigh_op_tnl_3')
// (16, 13, 'sp4_v_t_39')
// (16, 14, 'neigh_op_lft_3')
// (16, 14, 'sp4_v_b_39')
// (16, 15, 'neigh_op_bnl_3')
// (16, 15, 'sp4_v_b_26')
// (16, 16, 'sp4_v_b_15')
// (16, 17, 'sp4_v_b_2')
// (16, 17, 'sp4_v_t_39')
// (16, 18, 'sp4_v_b_39')
// (16, 19, 'sp4_v_b_26')
// (16, 20, 'local_g1_7')
// (16, 20, 'lutff_4/in_0')
// (16, 20, 'lutff_5/in_3')
// (16, 20, 'sp4_v_b_15')
// (16, 21, 'sp4_v_b_2')

reg n541 = 0;
// (11, 21, 'sp4_h_r_8')
// (12, 21, 'sp4_h_r_21')
// (13, 21, 'sp4_h_r_32')
// (14, 21, 'sp4_h_r_45')
// (14, 22, 'sp4_r_v_b_45')
// (14, 23, 'sp4_r_v_b_32')
// (14, 24, 'neigh_op_tnr_4')
// (14, 24, 'sp4_r_v_b_21')
// (14, 25, 'neigh_op_rgt_4')
// (14, 25, 'sp4_r_v_b_8')
// (14, 26, 'neigh_op_bnr_4')
// (15, 21, 'sp4_h_l_45')
// (15, 21, 'sp4_h_r_11')
// (15, 21, 'sp4_v_t_45')
// (15, 22, 'sp4_v_b_45')
// (15, 23, 'sp4_v_b_32')
// (15, 24, 'neigh_op_top_4')
// (15, 24, 'sp4_v_b_21')
// (15, 25, 'local_g3_4')
// (15, 25, 'lutff_4/in_1')
// (15, 25, 'lutff_4/out')
// (15, 25, 'sp4_v_b_8')
// (15, 26, 'neigh_op_bot_4')
// (16, 21, 'sp4_h_r_22')
// (16, 24, 'neigh_op_tnl_4')
// (16, 25, 'neigh_op_lft_4')
// (16, 26, 'neigh_op_bnl_4')
// (17, 21, 'sp4_h_r_35')
// (18, 21, 'local_g2_6')
// (18, 21, 'lutff_6/in_2')
// (18, 21, 'sp4_h_r_46')
// (19, 21, 'sp4_h_l_46')

wire n542;
// (11, 23, 'neigh_op_tnr_0')
// (11, 24, 'neigh_op_rgt_0')
// (11, 25, 'neigh_op_bnr_0')
// (12, 21, 'sp4_r_v_b_36')
// (12, 22, 'sp4_r_v_b_25')
// (12, 23, 'neigh_op_top_0')
// (12, 23, 'sp4_r_v_b_12')
// (12, 24, 'lutff_0/out')
// (12, 24, 'sp4_r_v_b_1')
// (12, 25, 'neigh_op_bot_0')
// (13, 20, 'sp4_v_t_36')
// (13, 21, 'local_g2_4')
// (13, 21, 'lutff_0/in_0')
// (13, 21, 'sp4_v_b_36')
// (13, 22, 'sp4_v_b_25')
// (13, 23, 'neigh_op_tnl_0')
// (13, 23, 'sp4_v_b_12')
// (13, 24, 'neigh_op_lft_0')
// (13, 24, 'sp4_v_b_1')
// (13, 25, 'neigh_op_bnl_0')

reg n543 = 0;
// (11, 24, 'sp12_h_r_1')
// (12, 24, 'sp12_h_r_2')
// (13, 24, 'sp12_h_r_5')
// (14, 24, 'sp12_h_r_6')
// (15, 23, 'neigh_op_tnr_1')
// (15, 24, 'neigh_op_rgt_1')
// (15, 24, 'sp12_h_r_9')
// (15, 25, 'neigh_op_bnr_1')
// (16, 23, 'neigh_op_top_1')
// (16, 24, 'lutff_1/out')
// (16, 24, 'sp12_h_r_10')
// (16, 25, 'neigh_op_bot_1')
// (17, 23, 'neigh_op_tnl_1')
// (17, 24, 'neigh_op_lft_1')
// (17, 24, 'sp12_h_r_13')
// (17, 25, 'neigh_op_bnl_1')
// (18, 24, 'sp12_h_r_14')
// (19, 24, 'sp12_h_r_17')
// (20, 24, 'sp12_h_r_18')
// (21, 24, 'sp12_h_r_21')
// (22, 24, 'sp12_h_r_22')
// (22, 28, 'sp4_r_v_b_42')
// (22, 29, 'sp4_r_v_b_31')
// (22, 30, 'sp4_r_v_b_18')
// (22, 31, 'sp4_r_v_b_7')
// (23, 24, 'sp12_h_l_22')
// (23, 24, 'sp12_v_t_22')
// (23, 25, 'sp12_v_b_22')
// (23, 26, 'sp12_v_b_21')
// (23, 27, 'sp12_v_b_18')
// (23, 27, 'sp4_v_t_42')
// (23, 28, 'sp12_v_b_17')
// (23, 28, 'sp4_v_b_42')
// (23, 29, 'sp12_v_b_14')
// (23, 29, 'sp4_v_b_31')
// (23, 30, 'sp12_v_b_13')
// (23, 30, 'sp4_v_b_18')
// (23, 31, 'sp12_v_b_10')
// (23, 31, 'sp4_h_r_1')
// (23, 31, 'sp4_v_b_7')
// (23, 32, 'sp12_v_b_9')
// (23, 33, 'span12_vert_6')
// (24, 31, 'sp4_h_r_12')
// (25, 31, 'sp4_h_r_25')
// (26, 31, 'sp4_h_r_36')
// (26, 32, 'sp4_r_v_b_36')
// (27, 31, 'sp4_h_l_36')
// (27, 31, 'sp4_v_t_36')
// (27, 32, 'sp4_v_b_36')
// (27, 33, 'span4_horz_r_0')
// (27, 33, 'span4_vert_25')
// (28, 33, 'span4_horz_r_4')
// (29, 33, 'span4_horz_r_8')
// (30, 33, 'io_0/D_OUT_0')
// (30, 33, 'local_g0_4')
// (30, 33, 'span4_horz_r_12')
// (31, 33, 'span4_horz_l_12')

wire n544;
// (12, 5, 'sp4_r_v_b_38')
// (12, 6, 'sp4_r_v_b_27')
// (12, 7, 'sp4_r_v_b_14')
// (12, 8, 'sp4_r_v_b_3')
// (13, 4, 'sp4_v_t_38')
// (13, 5, 'sp4_v_b_38')
// (13, 6, 'sp4_v_b_27')
// (13, 7, 'local_g0_6')
// (13, 7, 'lutff_3/in_1')
// (13, 7, 'sp4_v_b_14')
// (13, 8, 'sp4_h_r_10')
// (13, 8, 'sp4_v_b_3')
// (14, 7, 'neigh_op_tnr_1')
// (14, 8, 'neigh_op_rgt_1')
// (14, 8, 'sp4_h_r_23')
// (14, 9, 'neigh_op_bnr_1')
// (15, 7, 'neigh_op_top_1')
// (15, 8, 'lutff_1/out')
// (15, 8, 'sp4_h_r_34')
// (15, 9, 'neigh_op_bot_1')
// (16, 7, 'neigh_op_tnl_1')
// (16, 8, 'neigh_op_lft_1')
// (16, 8, 'sp4_h_r_47')
// (16, 9, 'neigh_op_bnl_1')
// (17, 8, 'sp4_h_l_47')

wire n545;
// (12, 7, 'neigh_op_tnr_6')
// (12, 8, 'neigh_op_rgt_6')
// (12, 8, 'sp4_h_r_1')
// (12, 9, 'neigh_op_bnr_6')
// (13, 7, 'neigh_op_top_6')
// (13, 8, 'lutff_6/out')
// (13, 8, 'sp4_h_r_12')
// (13, 9, 'neigh_op_bot_6')
// (14, 7, 'neigh_op_tnl_6')
// (14, 8, 'neigh_op_lft_6')
// (14, 8, 'sp4_h_r_25')
// (14, 9, 'neigh_op_bnl_6')
// (15, 8, 'local_g2_4')
// (15, 8, 'lutff_1/in_3')
// (15, 8, 'sp4_h_r_36')
// (16, 8, 'sp4_h_l_36')

reg n546 = 0;
// (12, 8, 'neigh_op_tnr_0')
// (12, 9, 'neigh_op_rgt_0')
// (12, 10, 'neigh_op_bnr_0')
// (13, 5, 'sp12_v_t_23')
// (13, 6, 'sp12_v_b_23')
// (13, 7, 'sp12_v_b_20')
// (13, 8, 'neigh_op_top_0')
// (13, 8, 'sp12_v_b_19')
// (13, 9, 'lutff_0/out')
// (13, 9, 'sp12_v_b_16')
// (13, 10, 'neigh_op_bot_0')
// (13, 10, 'sp12_v_b_15')
// (13, 11, 'sp12_v_b_12')
// (13, 12, 'sp12_v_b_11')
// (13, 13, 'local_g2_0')
// (13, 13, 'lutff_2/in_0')
// (13, 13, 'sp12_v_b_8')
// (13, 14, 'sp12_v_b_7')
// (13, 15, 'sp12_v_b_4')
// (13, 16, 'sp12_v_b_3')
// (13, 17, 'sp12_v_b_0')
// (14, 8, 'neigh_op_tnl_0')
// (14, 9, 'neigh_op_lft_0')
// (14, 10, 'neigh_op_bnl_0')

reg n547 = 0;
// (12, 8, 'neigh_op_tnr_2')
// (12, 9, 'neigh_op_rgt_2')
// (12, 9, 'sp4_r_v_b_36')
// (12, 10, 'neigh_op_bnr_2')
// (12, 10, 'sp4_r_v_b_25')
// (12, 11, 'sp4_r_v_b_12')
// (12, 12, 'sp4_r_v_b_1')
// (12, 13, 'sp4_r_v_b_41')
// (12, 14, 'sp4_r_v_b_28')
// (12, 15, 'sp4_r_v_b_17')
// (12, 16, 'sp4_r_v_b_4')
// (13, 8, 'neigh_op_top_2')
// (13, 8, 'sp4_v_t_36')
// (13, 9, 'lutff_2/out')
// (13, 9, 'sp4_v_b_36')
// (13, 10, 'neigh_op_bot_2')
// (13, 10, 'sp4_v_b_25')
// (13, 11, 'sp4_v_b_12')
// (13, 12, 'sp4_v_b_1')
// (13, 12, 'sp4_v_t_41')
// (13, 13, 'sp4_v_b_41')
// (13, 14, 'sp4_v_b_28')
// (13, 15, 'sp4_v_b_17')
// (13, 16, 'sp4_h_r_10')
// (13, 16, 'sp4_v_b_4')
// (14, 8, 'neigh_op_tnl_2')
// (14, 9, 'neigh_op_lft_2')
// (14, 10, 'neigh_op_bnl_2')
// (14, 16, 'local_g0_7')
// (14, 16, 'lutff_4/in_3')
// (14, 16, 'lutff_7/in_0')
// (14, 16, 'sp4_h_r_23')
// (15, 16, 'sp4_h_r_34')
// (16, 16, 'sp4_h_r_47')
// (17, 16, 'sp4_h_l_47')

reg n548 = 0;
// (12, 9, 'neigh_op_tnr_0')
// (12, 10, 'local_g3_0')
// (12, 10, 'lutff_7/in_0')
// (12, 10, 'neigh_op_rgt_0')
// (12, 11, 'neigh_op_bnr_0')
// (13, 9, 'neigh_op_top_0')
// (13, 10, 'lutff_0/out')
// (13, 11, 'neigh_op_bot_0')
// (14, 9, 'neigh_op_tnl_0')
// (14, 10, 'neigh_op_lft_0')
// (14, 11, 'neigh_op_bnl_0')

reg n549 = 0;
// (12, 9, 'neigh_op_tnr_1')
// (12, 10, 'neigh_op_rgt_1')
// (12, 11, 'neigh_op_bnr_1')
// (13, 8, 'sp4_r_v_b_43')
// (13, 9, 'neigh_op_top_1')
// (13, 9, 'sp4_r_v_b_30')
// (13, 10, 'lutff_1/out')
// (13, 10, 'sp4_r_v_b_19')
// (13, 11, 'neigh_op_bot_1')
// (13, 11, 'sp4_r_v_b_6')
// (13, 12, 'sp4_r_v_b_39')
// (13, 13, 'sp4_r_v_b_26')
// (13, 14, 'sp4_r_v_b_15')
// (13, 15, 'sp4_r_v_b_2')
// (14, 7, 'sp4_v_t_43')
// (14, 8, 'sp4_v_b_43')
// (14, 9, 'neigh_op_tnl_1')
// (14, 9, 'sp4_v_b_30')
// (14, 10, 'neigh_op_lft_1')
// (14, 10, 'sp4_v_b_19')
// (14, 11, 'neigh_op_bnl_1')
// (14, 11, 'sp4_v_b_6')
// (14, 11, 'sp4_v_t_39')
// (14, 12, 'local_g2_7')
// (14, 12, 'lutff_2/in_3')
// (14, 12, 'sp4_v_b_39')
// (14, 13, 'sp4_v_b_26')
// (14, 14, 'sp4_v_b_15')
// (14, 15, 'sp4_v_b_2')

reg n550 = 0;
// (12, 9, 'neigh_op_tnr_4')
// (12, 10, 'local_g3_4')
// (12, 10, 'lutff_1/in_0')
// (12, 10, 'neigh_op_rgt_4')
// (12, 11, 'neigh_op_bnr_4')
// (13, 9, 'neigh_op_top_4')
// (13, 10, 'lutff_4/out')
// (13, 11, 'neigh_op_bot_4')
// (14, 9, 'neigh_op_tnl_4')
// (14, 10, 'neigh_op_lft_4')
// (14, 11, 'neigh_op_bnl_4')

reg n551 = 0;
// (12, 9, 'neigh_op_tnr_7')
// (12, 10, 'local_g3_7')
// (12, 10, 'lutff_1/in_1')
// (12, 10, 'neigh_op_rgt_7')
// (12, 11, 'neigh_op_bnr_7')
// (13, 9, 'neigh_op_top_7')
// (13, 10, 'lutff_7/out')
// (13, 11, 'neigh_op_bot_7')
// (14, 9, 'neigh_op_tnl_7')
// (14, 10, 'neigh_op_lft_7')
// (14, 11, 'neigh_op_bnl_7')

reg n552 = 0;
// (12, 9, 'sp4_h_r_3')
// (13, 9, 'local_g1_6')
// (13, 9, 'lutff_2/in_3')
// (13, 9, 'sp4_h_r_14')
// (14, 8, 'neigh_op_tnr_3')
// (14, 9, 'neigh_op_rgt_3')
// (14, 9, 'sp4_h_r_27')
// (14, 10, 'neigh_op_bnr_3')
// (15, 8, 'neigh_op_top_3')
// (15, 9, 'lutff_3/out')
// (15, 9, 'sp4_h_r_38')
// (15, 10, 'neigh_op_bot_3')
// (16, 8, 'neigh_op_tnl_3')
// (16, 9, 'neigh_op_lft_3')
// (16, 9, 'sp4_h_l_38')
// (16, 10, 'neigh_op_bnl_3')

wire n553;
// (12, 9, 'sp4_r_v_b_37')
// (12, 10, 'local_g0_0')
// (12, 10, 'lutff_3/in_1')
// (12, 10, 'sp4_r_v_b_24')
// (12, 11, 'sp4_r_v_b_13')
// (12, 12, 'sp4_r_v_b_0')
// (13, 8, 'sp4_v_t_37')
// (13, 9, 'sp4_v_b_37')
// (13, 10, 'sp4_v_b_24')
// (13, 11, 'neigh_op_tnr_1')
// (13, 11, 'sp4_v_b_13')
// (13, 12, 'neigh_op_rgt_1')
// (13, 12, 'sp4_h_r_7')
// (13, 12, 'sp4_v_b_0')
// (13, 13, 'neigh_op_bnr_1')
// (14, 11, 'neigh_op_top_1')
// (14, 12, 'lutff_1/out')
// (14, 12, 'sp4_h_r_18')
// (14, 13, 'neigh_op_bot_1')
// (15, 11, 'neigh_op_tnl_1')
// (15, 12, 'neigh_op_lft_1')
// (15, 12, 'sp4_h_r_31')
// (15, 13, 'neigh_op_bnl_1')
// (16, 12, 'sp4_h_r_42')
// (17, 12, 'sp4_h_l_42')

reg n554 = 0;
// (12, 10, 'local_g1_1')
// (12, 10, 'lutff_7/in_1')
// (12, 10, 'sp4_h_r_1')
// (13, 10, 'sp4_h_r_12')
// (14, 9, 'neigh_op_tnr_2')
// (14, 10, 'neigh_op_rgt_2')
// (14, 10, 'sp4_h_r_25')
// (14, 11, 'neigh_op_bnr_2')
// (15, 9, 'neigh_op_top_2')
// (15, 10, 'lutff_2/out')
// (15, 10, 'sp4_h_r_36')
// (15, 11, 'neigh_op_bot_2')
// (16, 9, 'neigh_op_tnl_2')
// (16, 10, 'neigh_op_lft_2')
// (16, 10, 'sp4_h_l_36')
// (16, 11, 'neigh_op_bnl_2')

wire n555;
// (12, 10, 'lutff_1/lout')
// (12, 10, 'lutff_2/in_2')

wire n556;
// (12, 10, 'lutff_2/lout')
// (12, 10, 'lutff_3/in_2')

wire n557;
// (12, 10, 'neigh_op_tnr_0')
// (12, 11, 'neigh_op_rgt_0')
// (12, 12, 'neigh_op_bnr_0')
// (13, 7, 'sp12_v_t_23')
// (13, 8, 'sp12_v_b_23')
// (13, 9, 'sp12_v_b_20')
// (13, 10, 'neigh_op_top_0')
// (13, 10, 'sp12_v_b_19')
// (13, 11, 'local_g1_0')
// (13, 11, 'lutff_0/out')
// (13, 11, 'lutff_4/in_3')
// (13, 11, 'sp12_v_b_16')
// (13, 12, 'neigh_op_bot_0')
// (13, 12, 'sp12_v_b_15')
// (13, 13, 'local_g2_4')
// (13, 13, 'lutff_0/in_0')
// (13, 13, 'sp12_v_b_12')
// (13, 14, 'sp12_v_b_11')
// (13, 15, 'sp12_v_b_8')
// (13, 16, 'sp12_v_b_7')
// (13, 17, 'sp12_v_b_4')
// (13, 18, 'sp12_v_b_3')
// (13, 19, 'sp12_v_b_0')
// (14, 10, 'neigh_op_tnl_0')
// (14, 11, 'neigh_op_lft_0')
// (14, 12, 'neigh_op_bnl_0')

wire n558;
// (12, 10, 'neigh_op_tnr_1')
// (12, 11, 'neigh_op_rgt_1')
// (12, 12, 'neigh_op_bnr_1')
// (13, 10, 'neigh_op_top_1')
// (13, 11, 'local_g3_1')
// (13, 11, 'lutff_1/out')
// (13, 11, 'lutff_5/in_3')
// (13, 12, 'local_g1_1')
// (13, 12, 'lutff_0/in_2')
// (13, 12, 'neigh_op_bot_1')
// (14, 10, 'neigh_op_tnl_1')
// (14, 11, 'neigh_op_lft_1')
// (14, 12, 'neigh_op_bnl_1')

reg n559 = 0;
// (12, 10, 'neigh_op_tnr_2')
// (12, 11, 'neigh_op_rgt_2')
// (12, 11, 'sp4_r_v_b_36')
// (12, 12, 'neigh_op_bnr_2')
// (12, 12, 'sp4_r_v_b_25')
// (12, 13, 'sp4_r_v_b_12')
// (12, 14, 'sp4_r_v_b_1')
// (13, 10, 'neigh_op_top_2')
// (13, 10, 'sp4_v_t_36')
// (13, 11, 'local_g2_2')
// (13, 11, 'lutff_1/in_1')
// (13, 11, 'lutff_2/in_2')
// (13, 11, 'lutff_2/out')
// (13, 11, 'lutff_4/in_2')
// (13, 11, 'sp4_v_b_36')
// (13, 12, 'local_g1_2')
// (13, 12, 'lutff_2/in_1')
// (13, 12, 'neigh_op_bot_2')
// (13, 12, 'sp4_v_b_25')
// (13, 13, 'local_g1_4')
// (13, 13, 'lutff_0/in_1')
// (13, 13, 'sp4_v_b_12')
// (13, 14, 'sp4_v_b_1')
// (14, 10, 'neigh_op_tnl_2')
// (14, 11, 'neigh_op_lft_2')
// (14, 12, 'neigh_op_bnl_2')

reg n560 = 0;
// (12, 10, 'neigh_op_tnr_3')
// (12, 11, 'neigh_op_rgt_3')
// (12, 12, 'neigh_op_bnr_3')
// (13, 10, 'neigh_op_top_3')
// (13, 11, 'local_g0_3')
// (13, 11, 'lutff_0/in_1')
// (13, 11, 'lutff_3/in_0')
// (13, 11, 'lutff_3/out')
// (13, 12, 'local_g1_3')
// (13, 12, 'lutff_1/in_1')
// (13, 12, 'neigh_op_bot_3')
// (14, 10, 'neigh_op_tnl_3')
// (14, 11, 'neigh_op_lft_3')
// (14, 12, 'neigh_op_bnl_3')

wire n561;
// (12, 10, 'neigh_op_tnr_4')
// (12, 11, 'neigh_op_rgt_4')
// (12, 12, 'neigh_op_bnr_4')
// (13, 10, 'neigh_op_top_4')
// (13, 11, 'local_g0_4')
// (13, 11, 'lutff_2/in_0')
// (13, 11, 'lutff_3/in_1')
// (13, 11, 'lutff_4/out')
// (13, 12, 'neigh_op_bot_4')
// (14, 10, 'neigh_op_tnl_4')
// (14, 11, 'neigh_op_lft_4')
// (14, 12, 'neigh_op_bnl_4')

reg n562 = 0;
// (12, 10, 'neigh_op_tnr_5')
// (12, 11, 'neigh_op_rgt_5')
// (12, 12, 'neigh_op_bnr_5')
// (13, 10, 'neigh_op_top_5')
// (13, 11, 'local_g3_5')
// (13, 11, 'lutff_0/in_2')
// (13, 11, 'lutff_5/in_1')
// (13, 11, 'lutff_5/out')
// (13, 12, 'local_g0_5')
// (13, 12, 'lutff_0/in_1')
// (13, 12, 'neigh_op_bot_5')
// (14, 10, 'neigh_op_tnl_5')
// (14, 11, 'neigh_op_lft_5')
// (14, 12, 'neigh_op_bnl_5')

wire n563;
// (12, 10, 'neigh_op_tnr_6')
// (12, 10, 'sp4_r_v_b_41')
// (12, 11, 'neigh_op_rgt_6')
// (12, 11, 'sp4_r_v_b_28')
// (12, 11, 'sp4_r_v_b_44')
// (12, 12, 'local_g0_2')
// (12, 12, 'lutff_global/cen')
// (12, 12, 'neigh_op_bnr_6')
// (12, 12, 'sp4_r_v_b_17')
// (12, 12, 'sp4_r_v_b_33')
// (12, 13, 'sp4_r_v_b_20')
// (12, 13, 'sp4_r_v_b_4')
// (12, 14, 'sp4_r_v_b_9')
// (13, 9, 'sp4_v_t_41')
// (13, 10, 'neigh_op_top_6')
// (13, 10, 'sp4_v_b_41')
// (13, 10, 'sp4_v_t_44')
// (13, 11, 'lutff_6/out')
// (13, 11, 'sp4_v_b_28')
// (13, 11, 'sp4_v_b_44')
// (13, 12, 'neigh_op_bot_6')
// (13, 12, 'sp4_v_b_17')
// (13, 12, 'sp4_v_b_33')
// (13, 13, 'local_g0_2')
// (13, 13, 'lutff_global/cen')
// (13, 13, 'sp4_h_r_10')
// (13, 13, 'sp4_v_b_20')
// (13, 13, 'sp4_v_b_4')
// (13, 14, 'sp4_v_b_9')
// (14, 10, 'neigh_op_tnl_6')
// (14, 11, 'neigh_op_lft_6')
// (14, 12, 'neigh_op_bnl_6')
// (14, 13, 'sp4_h_r_23')
// (15, 13, 'sp4_h_r_34')
// (16, 13, 'sp4_h_r_47')
// (17, 13, 'sp4_h_l_47')

reg n564 = 0;
// (12, 10, 'sp12_h_r_1')
// (13, 10, 'sp12_h_r_2')
// (14, 10, 'local_g1_5')
// (14, 10, 'lutff_0/in_0')
// (14, 10, 'sp12_h_r_5')
// (15, 10, 'sp12_h_r_6')
// (16, 9, 'neigh_op_tnr_1')
// (16, 10, 'neigh_op_rgt_1')
// (16, 10, 'sp12_h_r_9')
// (16, 11, 'neigh_op_bnr_1')
// (17, 9, 'neigh_op_top_1')
// (17, 10, 'lutff_1/out')
// (17, 10, 'sp12_h_r_10')
// (17, 11, 'neigh_op_bot_1')
// (18, 9, 'neigh_op_tnl_1')
// (18, 10, 'neigh_op_lft_1')
// (18, 10, 'sp12_h_r_13')
// (18, 11, 'neigh_op_bnl_1')
// (19, 10, 'sp12_h_r_14')
// (20, 10, 'sp12_h_r_17')
// (21, 10, 'sp12_h_r_18')
// (22, 10, 'sp12_h_r_21')
// (23, 10, 'sp12_h_r_22')
// (24, 10, 'sp12_h_l_22')

wire n565;
// (12, 11, 'neigh_op_tnr_1')
// (12, 12, 'neigh_op_rgt_1')
// (12, 13, 'neigh_op_bnr_1')
// (13, 11, 'local_g1_1')
// (13, 11, 'lutff_3/in_3')
// (13, 11, 'neigh_op_top_1')
// (13, 12, 'lutff_1/out')
// (13, 13, 'neigh_op_bot_1')
// (14, 11, 'neigh_op_tnl_1')
// (14, 12, 'neigh_op_lft_1')
// (14, 13, 'neigh_op_bnl_1')

wire n566;
// (12, 11, 'neigh_op_tnr_2')
// (12, 12, 'neigh_op_rgt_2')
// (12, 13, 'neigh_op_bnr_2')
// (13, 11, 'local_g1_2')
// (13, 11, 'lutff_2/in_3')
// (13, 11, 'neigh_op_top_2')
// (13, 12, 'lutff_2/out')
// (13, 13, 'neigh_op_bot_2')
// (14, 11, 'neigh_op_tnl_2')
// (14, 12, 'neigh_op_lft_2')
// (14, 13, 'neigh_op_bnl_2')

reg n567 = 0;
// (12, 11, 'neigh_op_tnr_3')
// (12, 12, 'neigh_op_rgt_3')
// (12, 13, 'neigh_op_bnr_3')
// (13, 11, 'local_g1_3')
// (13, 11, 'lutff_0/in_0')
// (13, 11, 'neigh_op_top_3')
// (13, 12, 'local_g3_3')
// (13, 12, 'lutff_3/in_1')
// (13, 12, 'lutff_3/out')
// (13, 13, 'neigh_op_bot_3')
// (14, 11, 'neigh_op_tnl_3')
// (14, 12, 'neigh_op_lft_3')
// (14, 13, 'neigh_op_bnl_3')

reg n568 = 0;
// (12, 11, 'neigh_op_tnr_4')
// (12, 12, 'neigh_op_rgt_4')
// (12, 13, 'neigh_op_bnr_4')
// (13, 11, 'local_g1_4')
// (13, 11, 'lutff_0/in_3')
// (13, 11, 'neigh_op_top_4')
// (13, 12, 'local_g3_4')
// (13, 12, 'lutff_4/in_1')
// (13, 12, 'lutff_4/out')
// (13, 13, 'neigh_op_bot_4')
// (14, 11, 'neigh_op_tnl_4')
// (14, 12, 'neigh_op_lft_4')
// (14, 13, 'neigh_op_bnl_4')

reg n569 = 0;
// (12, 11, 'neigh_op_tnr_5')
// (12, 12, 'neigh_op_rgt_5')
// (12, 13, 'neigh_op_bnr_5')
// (13, 11, 'local_g1_5')
// (13, 11, 'lutff_1/in_3')
// (13, 11, 'lutff_4/in_0')
// (13, 11, 'neigh_op_top_5')
// (13, 12, 'local_g3_5')
// (13, 12, 'lutff_5/in_1')
// (13, 12, 'lutff_5/out')
// (13, 13, 'local_g0_5')
// (13, 13, 'lutff_0/in_3')
// (13, 13, 'neigh_op_bot_5')
// (14, 11, 'neigh_op_tnl_5')
// (14, 12, 'neigh_op_lft_5')
// (14, 13, 'neigh_op_bnl_5')

reg n570 = 0;
// (12, 11, 'sp12_h_r_1')
// (13, 11, 'sp12_h_r_2')
// (14, 11, 'sp12_h_r_5')
// (15, 11, 'sp12_h_r_6')
// (16, 11, 'sp12_h_r_9')
// (17, 11, 'local_g0_2')
// (17, 11, 'lutff_1/in_1')
// (17, 11, 'sp12_h_r_10')
// (18, 11, 'sp12_h_r_13')
// (19, 11, 'sp12_h_r_14')
// (20, 10, 'neigh_op_tnr_5')
// (20, 11, 'neigh_op_rgt_5')
// (20, 11, 'sp12_h_r_17')
// (20, 12, 'neigh_op_bnr_5')
// (21, 10, 'neigh_op_top_5')
// (21, 11, 'lutff_5/out')
// (21, 11, 'sp12_h_r_18')
// (21, 12, 'neigh_op_bot_5')
// (22, 10, 'neigh_op_tnl_5')
// (22, 11, 'neigh_op_lft_5')
// (22, 11, 'sp12_h_r_21')
// (22, 12, 'neigh_op_bnl_5')
// (23, 11, 'sp12_h_r_22')
// (24, 11, 'sp12_h_l_22')

reg n571 = 0;
// (12, 12, 'neigh_op_tnr_0')
// (12, 13, 'neigh_op_rgt_0')
// (12, 13, 'sp4_h_r_5')
// (12, 14, 'neigh_op_bnr_0')
// (13, 12, 'neigh_op_top_0')
// (13, 13, 'lutff_0/out')
// (13, 13, 'sp4_h_r_16')
// (13, 14, 'neigh_op_bot_0')
// (14, 12, 'neigh_op_tnl_0')
// (14, 13, 'neigh_op_lft_0')
// (14, 13, 'sp4_h_r_29')
// (14, 14, 'neigh_op_bnl_0')
// (15, 10, 'sp4_r_v_b_46')
// (15, 11, 'sp4_r_v_b_35')
// (15, 12, 'local_g3_6')
// (15, 12, 'lutff_5/in_0')
// (15, 12, 'sp4_r_v_b_22')
// (15, 13, 'sp4_h_r_40')
// (15, 13, 'sp4_r_v_b_11')
// (16, 9, 'sp4_v_t_46')
// (16, 10, 'sp4_v_b_46')
// (16, 11, 'sp4_v_b_35')
// (16, 12, 'sp4_v_b_22')
// (16, 13, 'sp4_h_l_40')
// (16, 13, 'sp4_v_b_11')

wire n572;
// (12, 12, 'neigh_op_tnr_3')
// (12, 13, 'neigh_op_rgt_3')
// (12, 14, 'local_g1_3')
// (12, 14, 'lutff_0/in_2')
// (12, 14, 'neigh_op_bnr_3')
// (13, 12, 'neigh_op_top_3')
// (13, 13, 'lutff_3/out')
// (13, 14, 'neigh_op_bot_3')
// (14, 12, 'neigh_op_tnl_3')
// (14, 13, 'neigh_op_lft_3')
// (14, 14, 'neigh_op_bnl_3')

wire n573;
// (12, 13, 'local_g1_3')
// (12, 13, 'lutff_global/cen')
// (12, 13, 'sp4_h_r_3')
// (13, 13, 'sp4_h_r_14')
// (14, 12, 'neigh_op_tnr_3')
// (14, 13, 'neigh_op_rgt_3')
// (14, 13, 'sp4_h_r_27')
// (14, 14, 'neigh_op_bnr_3')
// (15, 12, 'neigh_op_top_3')
// (15, 13, 'lutff_3/out')
// (15, 13, 'sp4_h_r_38')
// (15, 14, 'neigh_op_bot_3')
// (16, 12, 'neigh_op_tnl_3')
// (16, 13, 'neigh_op_lft_3')
// (16, 13, 'sp4_h_l_38')
// (16, 14, 'neigh_op_bnl_3')

reg n574 = 0;
// (12, 13, 'neigh_op_tnr_4')
// (12, 14, 'neigh_op_rgt_4')
// (12, 15, 'neigh_op_bnr_4')
// (13, 13, 'neigh_op_top_4')
// (13, 14, 'lutff_4/out')
// (13, 14, 'sp12_h_r_0')
// (13, 15, 'neigh_op_bot_4')
// (14, 13, 'neigh_op_tnl_4')
// (14, 14, 'neigh_op_lft_4')
// (14, 14, 'sp12_h_r_3')
// (14, 15, 'neigh_op_bnl_4')
// (15, 14, 'sp12_h_r_4')
// (16, 14, 'sp12_h_r_7')
// (17, 14, 'sp12_h_r_8')
// (18, 14, 'sp12_h_r_11')
// (18, 14, 'sp4_h_r_7')
// (19, 14, 'sp12_h_r_12')
// (19, 14, 'sp4_h_r_18')
// (20, 14, 'sp12_h_r_15')
// (20, 14, 'sp4_h_r_31')
// (21, 14, 'sp12_h_r_16')
// (21, 14, 'sp4_h_r_42')
// (21, 15, 'sp4_r_v_b_37')
// (21, 16, 'sp4_r_v_b_24')
// (21, 17, 'sp4_r_v_b_13')
// (21, 18, 'sp4_r_v_b_0')
// (22, 14, 'sp12_h_r_19')
// (22, 14, 'sp4_h_l_42')
// (22, 14, 'sp4_v_t_37')
// (22, 15, 'sp4_v_b_37')
// (22, 16, 'local_g2_0')
// (22, 16, 'lutff_1/in_1')
// (22, 16, 'sp4_v_b_24')
// (22, 17, 'sp4_v_b_13')
// (22, 18, 'sp4_v_b_0')
// (23, 14, 'sp12_h_r_20')
// (24, 14, 'sp12_h_r_23')
// (25, 14, 'sp12_h_l_23')

reg n575 = 0;
// (12, 13, 'sp12_h_r_1')
// (12, 25, 'sp12_h_r_1')
// (13, 13, 'sp12_h_r_2')
// (13, 25, 'sp12_h_r_2')
// (14, 13, 'sp12_h_r_5')
// (14, 25, 'sp12_h_r_5')
// (15, 13, 'sp12_h_r_6')
// (15, 25, 'sp12_h_r_6')
// (16, 10, 'sp4_r_v_b_40')
// (16, 11, 'sp4_r_v_b_29')
// (16, 12, 'sp4_r_v_b_16')
// (16, 13, 'sp12_h_r_9')
// (16, 13, 'sp4_r_v_b_5')
// (16, 14, 'sp4_r_v_b_40')
// (16, 15, 'sp4_r_v_b_29')
// (16, 16, 'sp4_r_v_b_16')
// (16, 17, 'sp4_r_v_b_5')
// (16, 18, 'sp4_r_v_b_40')
// (16, 19, 'sp4_r_v_b_29')
// (16, 20, 'sp4_r_v_b_16')
// (16, 21, 'sp4_r_v_b_5')
// (16, 22, 'sp4_r_v_b_39')
// (16, 23, 'sp4_r_v_b_26')
// (16, 24, 'neigh_op_tnr_1')
// (16, 24, 'sp4_r_v_b_15')
// (16, 25, 'neigh_op_rgt_1')
// (16, 25, 'sp12_h_r_9')
// (16, 25, 'sp4_h_r_7')
// (16, 25, 'sp4_r_v_b_2')
// (16, 26, 'neigh_op_bnr_1')
// (17, 9, 'sp4_v_t_40')
// (17, 10, 'local_g3_0')
// (17, 10, 'lutff_0/in_1')
// (17, 10, 'sp12_v_t_22')
// (17, 10, 'sp4_v_b_40')
// (17, 11, 'local_g3_5')
// (17, 11, 'local_g3_6')
// (17, 11, 'lutff_0/in_0')
// (17, 11, 'lutff_1/in_0')
// (17, 11, 'lutff_3/in_2')
// (17, 11, 'lutff_5/in_0')
// (17, 11, 'sp12_v_b_22')
// (17, 11, 'sp4_v_b_29')
// (17, 12, 'local_g2_5')
// (17, 12, 'local_g3_5')
// (17, 12, 'lutff_2/in_1')
// (17, 12, 'lutff_3/in_0')
// (17, 12, 'lutff_4/in_0')
// (17, 12, 'lutff_5/in_0')
// (17, 12, 'lutff_6/in_0')
// (17, 12, 'lutff_7/in_0')
// (17, 12, 'sp12_v_b_21')
// (17, 12, 'sp4_r_v_b_36')
// (17, 12, 'sp4_v_b_16')
// (17, 13, 'local_g2_2')
// (17, 13, 'local_g3_2')
// (17, 13, 'lutff_1/in_2')
// (17, 13, 'lutff_2/in_0')
// (17, 13, 'lutff_5/in_2')
// (17, 13, 'lutff_7/in_1')
// (17, 13, 'sp12_h_r_10')
// (17, 13, 'sp12_v_b_18')
// (17, 13, 'sp4_r_v_b_25')
// (17, 13, 'sp4_v_b_5')
// (17, 13, 'sp4_v_t_40')
// (17, 14, 'local_g3_0')
// (17, 14, 'local_g3_1')
// (17, 14, 'lutff_0/in_2')
// (17, 14, 'lutff_1/in_1')
// (17, 14, 'lutff_3/in_2')
// (17, 14, 'lutff_4/in_0')
// (17, 14, 'lutff_6/in_2')
// (17, 14, 'lutff_7/in_0')
// (17, 14, 'sp12_h_r_1')
// (17, 14, 'sp12_v_b_17')
// (17, 14, 'sp12_v_t_22')
// (17, 14, 'sp4_r_v_b_12')
// (17, 14, 'sp4_v_b_40')
// (17, 15, 'local_g2_5')
// (17, 15, 'local_g2_6')
// (17, 15, 'lutff_0/in_2')
// (17, 15, 'lutff_1/in_0')
// (17, 15, 'lutff_3/in_2')
// (17, 15, 'lutff_4/in_1')
// (17, 15, 'lutff_5/in_2')
// (17, 15, 'lutff_6/in_0')
// (17, 15, 'lutff_7/in_2')
// (17, 15, 'sp12_v_b_14')
// (17, 15, 'sp12_v_b_22')
// (17, 15, 'sp4_r_v_b_1')
// (17, 15, 'sp4_v_b_29')
// (17, 16, 'local_g3_5')
// (17, 16, 'lutff_0/in_2')
// (17, 16, 'lutff_2/in_2')
// (17, 16, 'lutff_3/in_1')
// (17, 16, 'lutff_4/in_2')
// (17, 16, 'sp12_v_b_13')
// (17, 16, 'sp12_v_b_21')
// (17, 16, 'sp4_r_v_b_42')
// (17, 16, 'sp4_r_v_b_47')
// (17, 16, 'sp4_v_b_16')
// (17, 17, 'local_g1_7')
// (17, 17, 'local_g3_2')
// (17, 17, 'lutff_0/in_2')
// (17, 17, 'lutff_1/in_0')
// (17, 17, 'lutff_3/in_0')
// (17, 17, 'lutff_7/in_0')
// (17, 17, 'sp12_v_b_10')
// (17, 17, 'sp12_v_b_18')
// (17, 17, 'sp4_r_v_b_31')
// (17, 17, 'sp4_r_v_b_34')
// (17, 17, 'sp4_v_b_5')
// (17, 17, 'sp4_v_t_40')
// (17, 18, 'sp12_v_b_17')
// (17, 18, 'sp12_v_b_9')
// (17, 18, 'sp4_r_v_b_18')
// (17, 18, 'sp4_r_v_b_23')
// (17, 18, 'sp4_v_b_40')
// (17, 19, 'sp12_v_b_14')
// (17, 19, 'sp12_v_b_6')
// (17, 19, 'sp4_r_v_b_10')
// (17, 19, 'sp4_r_v_b_7')
// (17, 19, 'sp4_v_b_29')
// (17, 20, 'sp12_v_b_13')
// (17, 20, 'sp12_v_b_5')
// (17, 20, 'sp4_r_v_b_36')
// (17, 20, 'sp4_r_v_b_46')
// (17, 20, 'sp4_v_b_16')
// (17, 21, 'local_g0_2')
// (17, 21, 'local_g3_2')
// (17, 21, 'lutff_5/in_0')
// (17, 21, 'lutff_6/in_0')
// (17, 21, 'sp12_v_b_10')
// (17, 21, 'sp12_v_b_2')
// (17, 21, 'sp4_h_r_2')
// (17, 21, 'sp4_r_v_b_25')
// (17, 21, 'sp4_r_v_b_35')
// (17, 21, 'sp4_v_b_5')
// (17, 21, 'sp4_v_t_39')
// (17, 22, 'sp12_h_r_1')
// (17, 22, 'sp12_v_b_1')
// (17, 22, 'sp12_v_b_9')
// (17, 22, 'sp12_v_t_22')
// (17, 22, 'sp4_r_v_b_12')
// (17, 22, 'sp4_r_v_b_22')
// (17, 22, 'sp4_v_b_39')
// (17, 23, 'sp12_v_b_22')
// (17, 23, 'sp12_v_b_6')
// (17, 23, 'sp4_r_v_b_1')
// (17, 23, 'sp4_r_v_b_11')
// (17, 23, 'sp4_v_b_26')
// (17, 24, 'neigh_op_top_1')
// (17, 24, 'sp12_v_b_21')
// (17, 24, 'sp12_v_b_5')
// (17, 24, 'sp4_r_v_b_46')
// (17, 24, 'sp4_v_b_15')
// (17, 25, 'local_g0_1')
// (17, 25, 'lutff_1/in_0')
// (17, 25, 'lutff_1/out')
// (17, 25, 'lutff_3/in_0')
// (17, 25, 'sp12_h_r_10')
// (17, 25, 'sp12_v_b_18')
// (17, 25, 'sp12_v_b_2')
// (17, 25, 'sp4_h_r_18')
// (17, 25, 'sp4_r_v_b_35')
// (17, 25, 'sp4_v_b_2')
// (17, 26, 'neigh_op_bot_1')
// (17, 26, 'sp12_v_b_1')
// (17, 26, 'sp12_v_b_17')
// (17, 26, 'sp4_r_v_b_22')
// (17, 27, 'sp12_v_b_14')
// (17, 27, 'sp4_r_v_b_11')
// (17, 28, 'sp12_v_b_13')
// (17, 29, 'sp12_v_b_10')
// (17, 30, 'sp12_v_b_9')
// (17, 31, 'sp12_v_b_6')
// (17, 32, 'sp12_v_b_5')
// (17, 33, 'span12_vert_2')
// (18, 11, 'sp4_v_t_36')
// (18, 12, 'sp4_v_b_36')
// (18, 13, 'sp12_h_r_13')
// (18, 13, 'sp4_v_b_25')
// (18, 14, 'sp12_h_r_2')
// (18, 14, 'sp4_v_b_12')
// (18, 15, 'local_g0_7')
// (18, 15, 'local_g1_1')
// (18, 15, 'lutff_2/in_2')
// (18, 15, 'lutff_3/in_0')
// (18, 15, 'lutff_5/in_1')
// (18, 15, 'sp4_h_r_7')
// (18, 15, 'sp4_v_b_1')
// (18, 15, 'sp4_v_t_42')
// (18, 15, 'sp4_v_t_47')
// (18, 16, 'local_g2_7')
// (18, 16, 'lutff_0/in_1')
// (18, 16, 'sp4_v_b_42')
// (18, 16, 'sp4_v_b_47')
// (18, 17, 'local_g2_7')
// (18, 17, 'local_g3_7')
// (18, 17, 'lutff_0/in_1')
// (18, 17, 'lutff_1/in_0')
// (18, 17, 'lutff_4/in_0')
// (18, 17, 'lutff_7/in_0')
// (18, 17, 'sp4_v_b_31')
// (18, 17, 'sp4_v_b_34')
// (18, 18, 'local_g1_2')
// (18, 18, 'local_g1_7')
// (18, 18, 'lutff_0/in_1')
// (18, 18, 'lutff_1/in_1')
// (18, 18, 'lutff_4/in_0')
// (18, 18, 'lutff_5/in_0')
// (18, 18, 'sp4_v_b_18')
// (18, 18, 'sp4_v_b_23')
// (18, 19, 'local_g0_7')
// (18, 19, 'local_g1_5')
// (18, 19, 'lutff_0/in_0')
// (18, 19, 'lutff_2/in_0')
// (18, 19, 'lutff_3/in_0')
// (18, 19, 'lutff_4/in_0')
// (18, 19, 'lutff_5/in_0')
// (18, 19, 'lutff_6/in_0')
// (18, 19, 'sp4_h_r_5')
// (18, 19, 'sp4_v_b_10')
// (18, 19, 'sp4_v_b_7')
// (18, 19, 'sp4_v_t_36')
// (18, 19, 'sp4_v_t_46')
// (18, 20, 'local_g2_4')
// (18, 20, 'local_g3_4')
// (18, 20, 'lutff_0/in_0')
// (18, 20, 'lutff_4/in_0')
// (18, 20, 'lutff_5/in_0')
// (18, 20, 'sp4_v_b_36')
// (18, 20, 'sp4_v_b_46')
// (18, 21, 'sp4_h_r_15')
// (18, 21, 'sp4_v_b_25')
// (18, 21, 'sp4_v_b_35')
// (18, 22, 'sp12_h_r_2')
// (18, 22, 'sp4_v_b_12')
// (18, 22, 'sp4_v_b_22')
// (18, 23, 'sp4_h_r_11')
// (18, 23, 'sp4_h_r_4')
// (18, 23, 'sp4_v_b_1')
// (18, 23, 'sp4_v_b_11')
// (18, 23, 'sp4_v_t_46')
// (18, 24, 'local_g3_1')
// (18, 24, 'local_g3_6')
// (18, 24, 'lutff_1/in_1')
// (18, 24, 'lutff_2/in_0')
// (18, 24, 'lutff_3/in_0')
// (18, 24, 'neigh_op_tnl_1')
// (18, 24, 'sp4_v_b_46')
// (18, 25, 'local_g2_7')
// (18, 25, 'local_g3_7')
// (18, 25, 'lutff_2/in_0')
// (18, 25, 'lutff_3/in_1')
// (18, 25, 'lutff_4/in_0')
// (18, 25, 'lutff_5/in_0')
// (18, 25, 'lutff_6/in_1')
// (18, 25, 'neigh_op_lft_1')
// (18, 25, 'sp12_h_r_13')
// (18, 25, 'sp4_h_r_31')
// (18, 25, 'sp4_v_b_35')
// (18, 26, 'local_g2_1')
// (18, 26, 'lutff_5/in_0')
// (18, 26, 'neigh_op_bnl_1')
// (18, 26, 'sp4_v_b_22')
// (18, 27, 'sp4_v_b_11')
// (19, 13, 'local_g0_6')
// (19, 13, 'local_g1_6')
// (19, 13, 'lutff_1/in_1')
// (19, 13, 'lutff_2/in_0')
// (19, 13, 'lutff_4/in_0')
// (19, 13, 'lutff_5/in_2')
// (19, 13, 'lutff_6/in_0')
// (19, 13, 'sp12_h_r_14')
// (19, 14, 'local_g3_0')
// (19, 14, 'local_g3_7')
// (19, 14, 'lutff_1/in_2')
// (19, 14, 'lutff_2/in_0')
// (19, 14, 'lutff_3/in_1')
// (19, 14, 'lutff_4/in_0')
// (19, 14, 'lutff_6/in_0')
// (19, 14, 'sp12_h_r_5')
// (19, 14, 'sp4_r_v_b_40')
// (19, 14, 'sp4_r_v_b_47')
// (19, 15, 'local_g0_5')
// (19, 15, 'lutff_2/in_1')
// (19, 15, 'lutff_4/in_1')
// (19, 15, 'lutff_7/in_0')
// (19, 15, 'sp4_h_r_18')
// (19, 15, 'sp4_r_v_b_29')
// (19, 15, 'sp4_r_v_b_34')
// (19, 16, 'sp4_r_v_b_16')
// (19, 16, 'sp4_r_v_b_23')
// (19, 17, 'sp4_r_v_b_10')
// (19, 17, 'sp4_r_v_b_5')
// (19, 18, 'local_g2_4')
// (19, 18, 'local_g3_2')
// (19, 18, 'lutff_1/in_2')
// (19, 18, 'lutff_2/in_0')
// (19, 18, 'lutff_3/in_2')
// (19, 18, 'lutff_4/in_0')
// (19, 18, 'lutff_6/in_0')
// (19, 18, 'sp4_r_v_b_36')
// (19, 18, 'sp4_r_v_b_42')
// (19, 18, 'sp4_r_v_b_44')
// (19, 19, 'sp4_h_r_16')
// (19, 19, 'sp4_r_v_b_25')
// (19, 19, 'sp4_r_v_b_31')
// (19, 19, 'sp4_r_v_b_33')
// (19, 20, 'sp4_r_v_b_12')
// (19, 20, 'sp4_r_v_b_18')
// (19, 20, 'sp4_r_v_b_20')
// (19, 21, 'sp4_h_r_26')
// (19, 21, 'sp4_r_v_b_1')
// (19, 21, 'sp4_r_v_b_7')
// (19, 21, 'sp4_r_v_b_9')
// (19, 22, 'sp12_h_r_5')
// (19, 22, 'sp4_r_v_b_36')
// (19, 22, 'sp4_r_v_b_42')
// (19, 23, 'sp4_h_r_17')
// (19, 23, 'sp4_h_r_22')
// (19, 23, 'sp4_r_v_b_25')
// (19, 23, 'sp4_r_v_b_31')
// (19, 24, 'sp4_r_v_b_12')
// (19, 24, 'sp4_r_v_b_18')
// (19, 25, 'sp12_h_r_14')
// (19, 25, 'sp4_h_r_42')
// (19, 25, 'sp4_r_v_b_1')
// (19, 25, 'sp4_r_v_b_7')
// (20, 13, 'local_g0_1')
// (20, 13, 'local_g1_1')
// (20, 13, 'lutff_0/in_0')
// (20, 13, 'lutff_1/in_0')
// (20, 13, 'lutff_3/in_0')
// (20, 13, 'lutff_6/in_0')
// (20, 13, 'sp12_h_r_17')
// (20, 13, 'sp4_v_t_40')
// (20, 13, 'sp4_v_t_47')
// (20, 14, 'sp12_h_r_6')
// (20, 14, 'sp4_v_b_40')
// (20, 14, 'sp4_v_b_47')
// (20, 15, 'sp4_h_r_31')
// (20, 15, 'sp4_v_b_29')
// (20, 15, 'sp4_v_b_34')
// (20, 16, 'sp4_v_b_16')
// (20, 16, 'sp4_v_b_23')
// (20, 17, 'local_g0_0')
// (20, 17, 'lutff_0/in_0')
// (20, 17, 'lutff_2/in_0')
// (20, 17, 'lutff_4/in_0')
// (20, 17, 'lutff_6/in_0')
// (20, 17, 'sp4_h_r_0')
// (20, 17, 'sp4_h_r_9')
// (20, 17, 'sp4_v_b_10')
// (20, 17, 'sp4_v_b_5')
// (20, 17, 'sp4_v_t_36')
// (20, 17, 'sp4_v_t_42')
// (20, 17, 'sp4_v_t_44')
// (20, 18, 'local_g2_4')
// (20, 18, 'lutff_0/in_0')
// (20, 18, 'lutff_5/in_1')
// (20, 18, 'sp4_v_b_36')
// (20, 18, 'sp4_v_b_42')
// (20, 18, 'sp4_v_b_44')
// (20, 19, 'sp4_h_r_29')
// (20, 19, 'sp4_v_b_25')
// (20, 19, 'sp4_v_b_31')
// (20, 19, 'sp4_v_b_33')
// (20, 20, 'sp4_v_b_12')
// (20, 20, 'sp4_v_b_18')
// (20, 20, 'sp4_v_b_20')
// (20, 21, 'local_g3_7')
// (20, 21, 'lutff_0/in_0')
// (20, 21, 'lutff_2/in_0')
// (20, 21, 'lutff_4/in_0')
// (20, 21, 'lutff_6/in_0')
// (20, 21, 'sp4_h_r_39')
// (20, 21, 'sp4_v_b_1')
// (20, 21, 'sp4_v_b_7')
// (20, 21, 'sp4_v_b_9')
// (20, 21, 'sp4_v_t_36')
// (20, 21, 'sp4_v_t_42')
// (20, 22, 'sp12_h_r_6')
// (20, 22, 'sp4_v_b_36')
// (20, 22, 'sp4_v_b_42')
// (20, 23, 'sp4_h_r_28')
// (20, 23, 'sp4_h_r_35')
// (20, 23, 'sp4_v_b_25')
// (20, 23, 'sp4_v_b_31')
// (20, 24, 'sp4_v_b_12')
// (20, 24, 'sp4_v_b_18')
// (20, 25, 'sp12_h_r_17')
// (20, 25, 'sp4_h_l_42')
// (20, 25, 'sp4_v_b_1')
// (20, 25, 'sp4_v_b_7')
// (21, 12, 'sp4_r_v_b_45')
// (21, 13, 'local_g1_2')
// (21, 13, 'local_g2_0')
// (21, 13, 'lutff_0/in_2')
// (21, 13, 'lutff_2/in_1')
// (21, 13, 'lutff_5/in_2')
// (21, 13, 'lutff_6/in_0')
// (21, 13, 'lutff_7/in_2')
// (21, 13, 'sp12_h_r_18')
// (21, 13, 'sp4_r_v_b_32')
// (21, 14, 'local_g0_1')
// (21, 14, 'local_g3_5')
// (21, 14, 'lutff_0/in_2')
// (21, 14, 'lutff_1/in_0')
// (21, 14, 'lutff_3/in_2')
// (21, 14, 'lutff_4/in_0')
// (21, 14, 'lutff_6/in_2')
// (21, 14, 'lutff_7/in_0')
// (21, 14, 'sp12_h_r_9')
// (21, 14, 'sp4_r_v_b_21')
// (21, 15, 'local_g2_2')
// (21, 15, 'local_g3_2')
// (21, 15, 'lutff_0/in_0')
// (21, 15, 'lutff_1/in_0')
// (21, 15, 'lutff_3/in_0')
// (21, 15, 'lutff_6/in_0')
// (21, 15, 'sp4_h_r_42')
// (21, 15, 'sp4_r_v_b_8')
// (21, 16, 'local_g3_0')
// (21, 16, 'local_g3_5')
// (21, 16, 'lutff_1/in_2')
// (21, 16, 'lutff_2/in_0')
// (21, 16, 'lutff_3/in_2')
// (21, 16, 'lutff_4/in_0')
// (21, 16, 'lutff_6/in_1')
// (21, 16, 'sp4_r_v_b_39')
// (21, 16, 'sp4_r_v_b_40')
// (21, 16, 'sp4_r_v_b_43')
// (21, 16, 'sp4_r_v_b_45')
// (21, 17, 'local_g0_6')
// (21, 17, 'lutff_0/in_0')
// (21, 17, 'lutff_2/in_0')
// (21, 17, 'lutff_4/in_2')
// (21, 17, 'lutff_6/in_0')
// (21, 17, 'sp4_h_r_13')
// (21, 17, 'sp4_h_r_20')
// (21, 17, 'sp4_r_v_b_26')
// (21, 17, 'sp4_r_v_b_29')
// (21, 17, 'sp4_r_v_b_30')
// (21, 17, 'sp4_r_v_b_32')
// (21, 18, 'local_g2_7')
// (21, 18, 'local_g3_5')
// (21, 18, 'lutff_0/in_3')
// (21, 18, 'lutff_1/in_0')
// (21, 18, 'lutff_3/in_2')
// (21, 18, 'lutff_4/in_0')
// (21, 18, 'lutff_6/in_3')
// (21, 18, 'lutff_7/in_1')
// (21, 18, 'sp4_r_v_b_15')
// (21, 18, 'sp4_r_v_b_16')
// (21, 18, 'sp4_r_v_b_19')
// (21, 18, 'sp4_r_v_b_21')
// (21, 19, 'sp4_h_r_40')
// (21, 19, 'sp4_r_v_b_2')
// (21, 19, 'sp4_r_v_b_5')
// (21, 19, 'sp4_r_v_b_6')
// (21, 19, 'sp4_r_v_b_8')
// (21, 20, 'sp4_r_v_b_40')
// (21, 20, 'sp4_r_v_b_46')
// (21, 20, 'sp4_r_v_b_47')
// (21, 21, 'local_g1_5')
// (21, 21, 'local_g2_3')
// (21, 21, 'lutff_0/in_0')
// (21, 21, 'lutff_4/in_2')
// (21, 21, 'lutff_5/in_0')
// (21, 21, 'sp4_h_l_39')
// (21, 21, 'sp4_r_v_b_29')
// (21, 21, 'sp4_r_v_b_34')
// (21, 21, 'sp4_r_v_b_35')
// (21, 22, 'local_g0_1')
// (21, 22, 'local_g3_7')
// (21, 22, 'lutff_0/in_0')
// (21, 22, 'lutff_1/in_0')
// (21, 22, 'lutff_2/in_0')
// (21, 22, 'lutff_3/in_0')
// (21, 22, 'lutff_5/in_0')
// (21, 22, 'sp12_h_r_9')
// (21, 22, 'sp4_r_v_b_16')
// (21, 22, 'sp4_r_v_b_22')
// (21, 22, 'sp4_r_v_b_23')
// (21, 23, 'sp4_h_r_41')
// (21, 23, 'sp4_h_r_46')
// (21, 23, 'sp4_r_v_b_10')
// (21, 23, 'sp4_r_v_b_11')
// (21, 23, 'sp4_r_v_b_5')
// (21, 25, 'sp12_h_r_18')
// (22, 11, 'sp4_v_t_45')
// (22, 12, 'sp4_v_b_45')
// (22, 13, 'local_g2_0')
// (22, 13, 'local_g3_0')
// (22, 13, 'lutff_0/in_2')
// (22, 13, 'lutff_1/in_1')
// (22, 13, 'lutff_3/in_2')
// (22, 13, 'lutff_4/in_0')
// (22, 13, 'lutff_6/in_2')
// (22, 13, 'lutff_7/in_0')
// (22, 13, 'sp12_h_r_21')
// (22, 13, 'sp4_v_b_32')
// (22, 14, 'sp12_h_r_10')
// (22, 14, 'sp4_v_b_21')
// (22, 15, 'sp4_h_l_42')
// (22, 15, 'sp4_v_b_8')
// (22, 15, 'sp4_v_t_39')
// (22, 15, 'sp4_v_t_40')
// (22, 15, 'sp4_v_t_43')
// (22, 15, 'sp4_v_t_45')
// (22, 16, 'local_g2_3')
// (22, 16, 'local_g3_7')
// (22, 16, 'lutff_1/in_2')
// (22, 16, 'lutff_2/in_0')
// (22, 16, 'lutff_4/in_1')
// (22, 16, 'lutff_5/in_2')
// (22, 16, 'lutff_6/in_0')
// (22, 16, 'sp4_v_b_39')
// (22, 16, 'sp4_v_b_40')
// (22, 16, 'sp4_v_b_43')
// (22, 16, 'sp4_v_b_45')
// (22, 17, 'sp4_h_r_24')
// (22, 17, 'sp4_h_r_33')
// (22, 17, 'sp4_v_b_26')
// (22, 17, 'sp4_v_b_29')
// (22, 17, 'sp4_v_b_30')
// (22, 17, 'sp4_v_b_32')
// (22, 18, 'sp4_v_b_15')
// (22, 18, 'sp4_v_b_16')
// (22, 18, 'sp4_v_b_19')
// (22, 18, 'sp4_v_b_21')
// (22, 19, 'local_g0_1')
// (22, 19, 'local_g1_5')
// (22, 19, 'lutff_2/in_1')
// (22, 19, 'lutff_4/in_0')
// (22, 19, 'lutff_6/in_0')
// (22, 19, 'lutff_7/in_0')
// (22, 19, 'sp4_h_l_40')
// (22, 19, 'sp4_h_r_1')
// (22, 19, 'sp4_v_b_2')
// (22, 19, 'sp4_v_b_5')
// (22, 19, 'sp4_v_b_6')
// (22, 19, 'sp4_v_b_8')
// (22, 19, 'sp4_v_t_40')
// (22, 19, 'sp4_v_t_46')
// (22, 19, 'sp4_v_t_47')
// (22, 20, 'local_g3_0')
// (22, 20, 'local_g3_7')
// (22, 20, 'lutff_1/in_0')
// (22, 20, 'lutff_2/in_0')
// (22, 20, 'lutff_6/in_0')
// (22, 20, 'lutff_7/in_0')
// (22, 20, 'sp4_v_b_40')
// (22, 20, 'sp4_v_b_46')
// (22, 20, 'sp4_v_b_47')
// (22, 21, 'sp4_v_b_29')
// (22, 21, 'sp4_v_b_34')
// (22, 21, 'sp4_v_b_35')
// (22, 22, 'sp12_h_r_10')
// (22, 22, 'sp4_v_b_16')
// (22, 22, 'sp4_v_b_22')
// (22, 22, 'sp4_v_b_23')
// (22, 23, 'sp4_h_l_41')
// (22, 23, 'sp4_h_l_46')
// (22, 23, 'sp4_v_b_10')
// (22, 23, 'sp4_v_b_11')
// (22, 23, 'sp4_v_b_5')
// (22, 25, 'sp12_h_r_21')
// (23, 13, 'local_g0_6')
// (23, 13, 'lutff_4/in_0')
// (23, 13, 'sp12_h_r_22')
// (23, 14, 'sp12_h_r_13')
// (23, 17, 'local_g3_4')
// (23, 17, 'lutff_2/in_1')
// (23, 17, 'lutff_4/in_1')
// (23, 17, 'lutff_7/in_0')
// (23, 17, 'sp4_h_r_37')
// (23, 17, 'sp4_h_r_44')
// (23, 19, 'local_g0_4')
// (23, 19, 'lutff_1/in_1')
// (23, 19, 'sp4_h_r_12')
// (23, 22, 'sp12_h_r_13')
// (23, 25, 'sp12_h_r_22')
// (24, 13, 'sp12_h_l_22')
// (24, 13, 'sp12_v_t_22')
// (24, 14, 'sp12_h_r_14')
// (24, 14, 'sp12_v_b_22')
// (24, 15, 'sp12_v_b_21')
// (24, 16, 'sp12_v_b_18')
// (24, 17, 'sp12_v_b_17')
// (24, 17, 'sp4_h_l_37')
// (24, 17, 'sp4_h_l_44')
// (24, 18, 'sp12_v_b_14')
// (24, 19, 'sp12_v_b_13')
// (24, 19, 'sp4_h_r_25')
// (24, 20, 'sp12_v_b_10')
// (24, 21, 'sp12_v_b_9')
// (24, 22, 'sp12_h_r_14')
// (24, 22, 'sp12_v_b_6')
// (24, 23, 'sp12_v_b_5')
// (24, 24, 'sp12_v_b_2')
// (24, 25, 'sp12_h_l_22')
// (24, 25, 'sp12_v_b_1')
// (25, 14, 'sp12_h_r_17')
// (25, 19, 'sp4_h_r_36')
// (25, 22, 'sp12_h_r_17')
// (26, 14, 'sp12_h_r_18')
// (26, 19, 'sp4_h_l_36')
// (26, 22, 'sp12_h_r_18')
// (27, 14, 'sp12_h_r_21')
// (27, 22, 'sp12_h_r_21')
// (28, 14, 'sp12_h_r_22')
// (28, 22, 'sp12_h_r_22')
// (29, 14, 'sp12_h_l_22')
// (29, 22, 'sp12_h_l_22')

wire n576;
// (12, 14, 'lutff_7/cout')
// (12, 15, 'carry_in')
// (12, 15, 'carry_in_mux')

reg n577 = 0;
// (12, 14, 'neigh_op_tnr_0')
// (12, 15, 'neigh_op_rgt_0')
// (12, 16, 'neigh_op_bnr_0')
// (13, 14, 'neigh_op_top_0')
// (13, 15, 'local_g2_0')
// (13, 15, 'lutff_0/out')
// (13, 15, 'lutff_1/in_3')
// (13, 16, 'neigh_op_bot_0')
// (14, 14, 'neigh_op_tnl_0')
// (14, 15, 'local_g0_0')
// (14, 15, 'lutff_5/in_1')
// (14, 15, 'neigh_op_lft_0')
// (14, 16, 'neigh_op_bnl_0')

reg n578 = 0;
// (12, 14, 'neigh_op_tnr_1')
// (12, 15, 'neigh_op_rgt_1')
// (12, 16, 'neigh_op_bnr_1')
// (13, 14, 'neigh_op_top_1')
// (13, 15, 'lutff_1/out')
// (13, 16, 'neigh_op_bot_1')
// (14, 14, 'neigh_op_tnl_1')
// (14, 15, 'local_g0_1')
// (14, 15, 'lutff_5/in_2')
// (14, 15, 'neigh_op_lft_1')
// (14, 16, 'neigh_op_bnl_1')

reg n579 = 0;
// (12, 14, 'neigh_op_tnr_2')
// (12, 15, 'neigh_op_rgt_2')
// (12, 16, 'neigh_op_bnr_2')
// (13, 14, 'neigh_op_top_2')
// (13, 15, 'local_g3_2')
// (13, 15, 'lutff_0/in_3')
// (13, 15, 'lutff_2/out')
// (13, 16, 'neigh_op_bot_2')
// (14, 14, 'neigh_op_tnl_2')
// (14, 15, 'local_g1_2')
// (14, 15, 'lutff_5/in_0')
// (14, 15, 'neigh_op_lft_2')
// (14, 16, 'neigh_op_bnl_2')

wire n580;
// (12, 14, 'sp4_h_r_7')
// (13, 14, 'local_g0_2')
// (13, 14, 'lutff_global/cen')
// (13, 14, 'sp4_h_r_18')
// (14, 14, 'sp4_h_r_31')
// (15, 13, 'neigh_op_tnr_2')
// (15, 14, 'neigh_op_rgt_2')
// (15, 14, 'sp4_h_r_42')
// (15, 15, 'neigh_op_bnr_2')
// (16, 13, 'neigh_op_top_2')
// (16, 14, 'lutff_2/out')
// (16, 14, 'sp4_h_l_42')
// (16, 14, 'sp4_h_r_4')
// (16, 15, 'neigh_op_bot_2')
// (17, 13, 'neigh_op_tnl_2')
// (17, 14, 'neigh_op_lft_2')
// (17, 14, 'sp4_h_r_17')
// (17, 15, 'neigh_op_bnl_2')
// (18, 14, 'sp4_h_r_28')
// (19, 7, 'sp4_r_v_b_47')
// (19, 8, 'sp4_r_v_b_34')
// (19, 9, 'sp4_r_v_b_23')
// (19, 10, 'local_g2_2')
// (19, 10, 'lutff_global/cen')
// (19, 10, 'sp4_r_v_b_10')
// (19, 11, 'sp4_r_v_b_47')
// (19, 12, 'sp4_r_v_b_34')
// (19, 13, 'sp4_r_v_b_23')
// (19, 14, 'sp4_h_r_41')
// (19, 14, 'sp4_r_v_b_10')
// (20, 6, 'sp4_v_t_47')
// (20, 7, 'sp4_v_b_47')
// (20, 8, 'sp4_v_b_34')
// (20, 9, 'sp4_v_b_23')
// (20, 10, 'sp4_v_b_10')
// (20, 10, 'sp4_v_t_47')
// (20, 11, 'sp4_v_b_47')
// (20, 12, 'sp4_v_b_34')
// (20, 13, 'sp4_v_b_23')
// (20, 14, 'sp4_h_l_41')
// (20, 14, 'sp4_v_b_10')

wire n581;
// (12, 15, 'lutff_7/cout')
// (12, 16, 'carry_in')
// (12, 16, 'carry_in_mux')
// (12, 16, 'lutff_0/in_3')

reg n582 = 0;
// (12, 15, 'neigh_op_tnr_0')
// (12, 16, 'neigh_op_rgt_0')
// (12, 17, 'neigh_op_bnr_0')
// (13, 12, 'sp12_v_t_23')
// (13, 13, 'sp12_v_b_23')
// (13, 14, 'sp12_v_b_20')
// (13, 15, 'neigh_op_top_0')
// (13, 15, 'sp12_v_b_19')
// (13, 16, 'lutff_0/out')
// (13, 16, 'sp12_v_b_16')
// (13, 17, 'neigh_op_bot_0')
// (13, 17, 'sp12_v_b_15')
// (13, 18, 'sp12_v_b_12')
// (13, 19, 'local_g2_3')
// (13, 19, 'lutff_2/in_1')
// (13, 19, 'sp12_v_b_11')
// (13, 20, 'sp12_v_b_8')
// (13, 21, 'sp12_v_b_7')
// (13, 22, 'sp12_v_b_4')
// (13, 23, 'sp12_v_b_3')
// (13, 24, 'sp12_v_b_0')
// (14, 15, 'neigh_op_tnl_0')
// (14, 16, 'neigh_op_lft_0')
// (14, 17, 'neigh_op_bnl_0')

reg n583 = 0;
// (12, 15, 'neigh_op_tnr_1')
// (12, 16, 'neigh_op_rgt_1')
// (12, 17, 'neigh_op_bnr_1')
// (13, 13, 'sp12_v_t_22')
// (13, 14, 'sp12_v_b_22')
// (13, 15, 'neigh_op_top_1')
// (13, 15, 'sp12_v_b_21')
// (13, 16, 'lutff_1/out')
// (13, 16, 'sp12_v_b_18')
// (13, 17, 'neigh_op_bot_1')
// (13, 17, 'sp12_v_b_17')
// (13, 18, 'sp12_v_b_14')
// (13, 19, 'local_g2_5')
// (13, 19, 'lutff_3/in_2')
// (13, 19, 'sp12_v_b_13')
// (13, 20, 'sp12_v_b_10')
// (13, 21, 'sp12_v_b_9')
// (13, 22, 'sp12_v_b_6')
// (13, 23, 'sp12_v_b_5')
// (13, 24, 'sp12_v_b_2')
// (13, 25, 'sp12_v_b_1')
// (14, 15, 'neigh_op_tnl_1')
// (14, 16, 'neigh_op_lft_1')
// (14, 17, 'neigh_op_bnl_1')

reg n584 = 0;
// (12, 15, 'neigh_op_tnr_2')
// (12, 16, 'neigh_op_rgt_2')
// (12, 16, 'sp4_r_v_b_36')
// (12, 17, 'neigh_op_bnr_2')
// (12, 17, 'sp4_r_v_b_25')
// (12, 18, 'sp4_r_v_b_12')
// (12, 19, 'sp4_r_v_b_1')
// (13, 15, 'neigh_op_top_2')
// (13, 15, 'sp4_v_t_36')
// (13, 16, 'lutff_2/out')
// (13, 16, 'sp4_v_b_36')
// (13, 17, 'neigh_op_bot_2')
// (13, 17, 'sp4_v_b_25')
// (13, 18, 'sp4_v_b_12')
// (13, 19, 'local_g0_1')
// (13, 19, 'lutff_4/in_1')
// (13, 19, 'sp4_v_b_1')
// (14, 15, 'neigh_op_tnl_2')
// (14, 16, 'neigh_op_lft_2')
// (14, 17, 'neigh_op_bnl_2')

reg n585 = 0;
// (12, 15, 'neigh_op_tnr_3')
// (12, 16, 'neigh_op_rgt_3')
// (12, 17, 'neigh_op_bnr_3')
// (13, 15, 'neigh_op_top_3')
// (13, 15, 'sp12_v_t_22')
// (13, 16, 'lutff_3/out')
// (13, 16, 'sp12_v_b_22')
// (13, 17, 'neigh_op_bot_3')
// (13, 17, 'sp12_v_b_21')
// (13, 18, 'sp12_v_b_18')
// (13, 19, 'local_g2_1')
// (13, 19, 'lutff_5/in_2')
// (13, 19, 'sp12_v_b_17')
// (13, 20, 'sp12_v_b_14')
// (13, 21, 'sp12_v_b_13')
// (13, 22, 'sp12_v_b_10')
// (13, 23, 'sp12_v_b_9')
// (13, 24, 'sp12_v_b_6')
// (13, 25, 'sp12_v_b_5')
// (13, 26, 'sp12_v_b_2')
// (13, 27, 'sp12_v_b_1')
// (14, 15, 'neigh_op_tnl_3')
// (14, 16, 'neigh_op_lft_3')
// (14, 17, 'neigh_op_bnl_3')

reg n586 = 0;
// (12, 15, 'neigh_op_tnr_4')
// (12, 16, 'neigh_op_rgt_4')
// (12, 16, 'sp4_r_v_b_40')
// (12, 17, 'neigh_op_bnr_4')
// (12, 17, 'sp4_r_v_b_29')
// (12, 18, 'sp4_r_v_b_16')
// (12, 19, 'sp4_r_v_b_5')
// (13, 15, 'neigh_op_top_4')
// (13, 15, 'sp4_v_t_40')
// (13, 16, 'lutff_4/out')
// (13, 16, 'sp4_v_b_40')
// (13, 17, 'neigh_op_bot_4')
// (13, 17, 'sp4_v_b_29')
// (13, 18, 'sp4_v_b_16')
// (13, 19, 'local_g0_5')
// (13, 19, 'lutff_6/in_1')
// (13, 19, 'sp4_v_b_5')
// (14, 15, 'neigh_op_tnl_4')
// (14, 16, 'neigh_op_lft_4')
// (14, 17, 'neigh_op_bnl_4')

reg n587 = 0;
// (12, 15, 'neigh_op_tnr_5')
// (12, 16, 'neigh_op_rgt_5')
// (12, 16, 'sp4_r_v_b_42')
// (12, 17, 'neigh_op_bnr_5')
// (12, 17, 'sp4_r_v_b_31')
// (12, 18, 'sp4_r_v_b_18')
// (12, 19, 'sp4_r_v_b_7')
// (13, 15, 'neigh_op_top_5')
// (13, 15, 'sp4_v_t_42')
// (13, 16, 'lutff_5/out')
// (13, 16, 'sp4_v_b_42')
// (13, 17, 'neigh_op_bot_5')
// (13, 17, 'sp4_v_b_31')
// (13, 18, 'sp4_v_b_18')
// (13, 19, 'local_g0_7')
// (13, 19, 'lutff_7/in_2')
// (13, 19, 'sp4_v_b_7')
// (14, 15, 'neigh_op_tnl_5')
// (14, 16, 'neigh_op_lft_5')
// (14, 17, 'neigh_op_bnl_5')

reg n588 = 0;
// (12, 15, 'neigh_op_tnr_6')
// (12, 16, 'neigh_op_rgt_6')
// (12, 17, 'neigh_op_bnr_6')
// (13, 10, 'sp12_v_t_23')
// (13, 11, 'sp12_v_b_23')
// (13, 12, 'sp12_v_b_20')
// (13, 13, 'sp12_v_b_19')
// (13, 14, 'sp12_v_b_16')
// (13, 15, 'neigh_op_top_6')
// (13, 15, 'sp12_v_b_15')
// (13, 16, 'lutff_6/out')
// (13, 16, 'sp12_v_b_12')
// (13, 17, 'neigh_op_bot_6')
// (13, 17, 'sp12_v_b_11')
// (13, 18, 'sp12_v_b_8')
// (13, 19, 'local_g2_7')
// (13, 19, 'lutff_0/in_1')
// (13, 19, 'sp12_v_b_7')
// (13, 20, 'sp12_v_b_4')
// (13, 21, 'sp12_v_b_3')
// (13, 22, 'sp12_v_b_0')
// (14, 15, 'neigh_op_tnl_6')
// (14, 16, 'neigh_op_lft_6')
// (14, 17, 'neigh_op_bnl_6')

reg n589 = 0;
// (12, 15, 'neigh_op_tnr_7')
// (12, 16, 'neigh_op_rgt_7')
// (12, 16, 'sp4_r_v_b_46')
// (12, 17, 'neigh_op_bnr_7')
// (12, 17, 'sp4_r_v_b_35')
// (12, 18, 'sp4_r_v_b_22')
// (12, 19, 'sp4_r_v_b_11')
// (13, 15, 'neigh_op_top_7')
// (13, 15, 'sp4_v_t_46')
// (13, 16, 'lutff_7/out')
// (13, 16, 'sp4_v_b_46')
// (13, 17, 'neigh_op_bot_7')
// (13, 17, 'sp4_v_b_35')
// (13, 18, 'sp4_v_b_22')
// (13, 19, 'local_g0_3')
// (13, 19, 'lutff_1/in_2')
// (13, 19, 'sp4_v_b_11')
// (14, 15, 'neigh_op_tnl_7')
// (14, 16, 'neigh_op_lft_7')
// (14, 17, 'neigh_op_bnl_7')

wire n590;
// (12, 15, 'sp12_h_r_0')
// (13, 15, 'sp12_h_r_3')
// (14, 15, 'sp12_h_r_4')
// (15, 13, 'sp4_r_v_b_40')
// (15, 14, 'neigh_op_tnr_0')
// (15, 14, 'sp4_r_v_b_29')
// (15, 15, 'neigh_op_rgt_0')
// (15, 15, 'sp12_h_r_7')
// (15, 15, 'sp4_r_v_b_16')
// (15, 16, 'local_g1_0')
// (15, 16, 'lutff_2/in_3')
// (15, 16, 'neigh_op_bnr_0')
// (15, 16, 'sp4_r_v_b_5')
// (15, 17, 'sp4_r_v_b_40')
// (15, 18, 'sp4_r_v_b_29')
// (15, 19, 'sp4_r_v_b_16')
// (15, 20, 'sp4_r_v_b_5')
// (16, 12, 'sp4_h_r_10')
// (16, 12, 'sp4_v_t_40')
// (16, 13, 'local_g3_0')
// (16, 13, 'lutff_0/in_3')
// (16, 13, 'lutff_5/in_0')
// (16, 13, 'lutff_7/in_0')
// (16, 13, 'sp4_v_b_40')
// (16, 14, 'neigh_op_top_0')
// (16, 14, 'sp4_v_b_29')
// (16, 15, 'lutff_0/out')
// (16, 15, 'sp12_h_r_8')
// (16, 15, 'sp4_v_b_16')
// (16, 16, 'neigh_op_bot_0')
// (16, 16, 'sp4_v_b_5')
// (16, 16, 'sp4_v_t_40')
// (16, 17, 'sp4_v_b_40')
// (16, 18, 'sp4_v_b_29')
// (16, 19, 'sp4_v_b_16')
// (16, 20, 'sp4_h_r_11')
// (16, 20, 'sp4_v_b_5')
// (17, 12, 'sp4_h_r_23')
// (17, 14, 'neigh_op_tnl_0')
// (17, 15, 'neigh_op_lft_0')
// (17, 15, 'sp12_h_r_11')
// (17, 16, 'neigh_op_bnl_0')
// (17, 20, 'sp4_h_r_22')
// (18, 12, 'sp4_h_r_34')
// (18, 15, 'sp12_h_r_12')
// (18, 20, 'sp4_h_r_35')
// (19, 12, 'local_g3_7')
// (19, 12, 'lutff_1/in_3')
// (19, 12, 'lutff_2/in_0')
// (19, 12, 'lutff_3/in_3')
// (19, 12, 'sp4_h_r_47')
// (19, 15, 'sp12_h_r_15')
// (19, 20, 'local_g3_6')
// (19, 20, 'lutff_6/in_3')
// (19, 20, 'lutff_7/in_0')
// (19, 20, 'sp4_h_r_46')
// (20, 12, 'sp4_h_l_47')
// (20, 15, 'local_g0_0')
// (20, 15, 'lutff_6/in_0')
// (20, 15, 'lutff_7/in_1')
// (20, 15, 'sp12_h_r_16')
// (20, 20, 'sp4_h_l_46')
// (21, 15, 'sp12_h_r_19')
// (22, 15, 'local_g1_4')
// (22, 15, 'lutff_0/in_3')
// (22, 15, 'lutff_4/in_3')
// (22, 15, 'lutff_5/in_0')
// (22, 15, 'sp12_h_r_20')
// (23, 15, 'sp12_h_r_23')
// (24, 15, 'sp12_h_l_23')

wire n591;
// (12, 15, 'sp4_h_r_2')
// (13, 12, 'sp4_r_v_b_47')
// (13, 13, 'sp4_r_v_b_34')
// (13, 14, 'neigh_op_tnr_5')
// (13, 14, 'sp4_r_v_b_23')
// (13, 15, 'neigh_op_rgt_5')
// (13, 15, 'sp4_h_r_15')
// (13, 15, 'sp4_r_v_b_10')
// (13, 16, 'neigh_op_bnr_5')
// (14, 11, 'sp4_v_t_47')
// (14, 12, 'local_g3_7')
// (14, 12, 'lutff_4/in_0')
// (14, 12, 'sp4_r_v_b_46')
// (14, 12, 'sp4_v_b_47')
// (14, 13, 'sp4_r_v_b_35')
// (14, 13, 'sp4_v_b_34')
// (14, 14, 'neigh_op_top_5')
// (14, 14, 'sp4_r_v_b_22')
// (14, 14, 'sp4_v_b_23')
// (14, 15, 'lutff_5/out')
// (14, 15, 'sp4_h_r_26')
// (14, 15, 'sp4_r_v_b_11')
// (14, 15, 'sp4_v_b_10')
// (14, 16, 'neigh_op_bot_5')
// (15, 11, 'sp4_v_t_46')
// (15, 12, 'local_g2_6')
// (15, 12, 'lutff_1/in_1')
// (15, 12, 'sp4_r_v_b_45')
// (15, 12, 'sp4_v_b_46')
// (15, 13, 'local_g3_3')
// (15, 13, 'lutff_2/in_0')
// (15, 13, 'lutff_3/in_3')
// (15, 13, 'sp4_r_v_b_32')
// (15, 13, 'sp4_v_b_35')
// (15, 14, 'local_g3_5')
// (15, 14, 'lutff_0/in_0')
// (15, 14, 'lutff_3/in_3')
// (15, 14, 'lutff_4/in_0')
// (15, 14, 'lutff_5/in_3')
// (15, 14, 'lutff_7/in_3')
// (15, 14, 'neigh_op_tnl_5')
// (15, 14, 'sp4_r_v_b_21')
// (15, 14, 'sp4_v_b_22')
// (15, 15, 'neigh_op_lft_5')
// (15, 15, 'sp4_h_r_39')
// (15, 15, 'sp4_r_v_b_8')
// (15, 15, 'sp4_v_b_11')
// (15, 16, 'neigh_op_bnl_5')
// (16, 11, 'sp4_v_t_45')
// (16, 12, 'local_g2_5')
// (16, 12, 'lutff_4/in_3')
// (16, 12, 'sp4_v_b_45')
// (16, 13, 'sp4_v_b_32')
// (16, 14, 'sp4_v_b_21')
// (16, 15, 'sp4_h_l_39')
// (16, 15, 'sp4_v_b_8')

wire n592;
// (12, 15, 'sp4_h_r_7')
// (13, 15, 'sp4_h_r_18')
// (14, 15, 'sp4_h_r_31')
// (15, 12, 'local_g2_4')
// (15, 12, 'lutff_0/in_0')
// (15, 12, 'sp4_r_v_b_36')
// (15, 13, 'sp4_r_v_b_25')
// (15, 14, 'sp4_r_v_b_12')
// (15, 15, 'sp4_h_r_42')
// (15, 15, 'sp4_r_v_b_1')
// (16, 11, 'sp4_v_t_36')
// (16, 12, 'sp4_v_b_36')
// (16, 13, 'sp4_v_b_25')
// (16, 14, 'sp4_v_b_12')
// (16, 15, 'sp4_h_l_42')
// (16, 15, 'sp4_h_r_11')
// (16, 15, 'sp4_v_b_1')
// (17, 15, 'sp4_h_r_22')
// (18, 15, 'sp4_h_r_35')
// (19, 14, 'neigh_op_tnr_4')
// (19, 15, 'neigh_op_rgt_4')
// (19, 15, 'sp4_h_r_46')
// (19, 16, 'neigh_op_bnr_4')
// (20, 14, 'neigh_op_top_4')
// (20, 15, 'local_g0_4')
// (20, 15, 'lutff_4/out')
// (20, 15, 'lutff_7/in_3')
// (20, 15, 'sp4_h_l_46')
// (20, 15, 'sp4_h_r_8')
// (20, 16, 'neigh_op_bot_4')
// (21, 14, 'neigh_op_tnl_4')
// (21, 15, 'neigh_op_lft_4')
// (21, 15, 'sp4_h_r_21')
// (21, 16, 'neigh_op_bnl_4')
// (22, 15, 'sp4_h_r_32')
// (23, 15, 'sp4_h_r_45')
// (24, 15, 'sp4_h_l_45')

wire n593;
// (12, 16, 'neigh_op_tnr_1')
// (12, 17, 'neigh_op_rgt_1')
// (12, 18, 'neigh_op_bnr_1')
// (13, 16, 'neigh_op_top_1')
// (13, 17, 'local_g0_1')
// (13, 17, 'lutff_1/out')
// (13, 17, 'lutff_4/in_1')
// (13, 18, 'neigh_op_bot_1')
// (14, 16, 'neigh_op_tnl_1')
// (14, 17, 'neigh_op_lft_1')
// (14, 18, 'neigh_op_bnl_1')

wire n594;
// (12, 16, 'neigh_op_tnr_7')
// (12, 17, 'neigh_op_rgt_7')
// (12, 18, 'neigh_op_bnr_7')
// (13, 16, 'neigh_op_top_7')
// (13, 17, 'local_g0_7')
// (13, 17, 'lutff_4/in_3')
// (13, 17, 'lutff_7/out')
// (13, 18, 'neigh_op_bot_7')
// (14, 16, 'neigh_op_tnl_7')
// (14, 17, 'neigh_op_lft_7')
// (14, 18, 'neigh_op_bnl_7')

reg n595 = 0;
// (12, 16, 'sp12_h_r_0')
// (13, 16, 'sp12_h_r_3')
// (14, 16, 'sp12_h_r_4')
// (14, 17, 'local_g0_1')
// (14, 17, 'lutff_3/in_0')
// (14, 17, 'sp4_h_r_9')
// (15, 16, 'sp12_h_r_7')
// (15, 17, 'sp4_h_r_20')
// (16, 16, 'sp12_h_r_8')
// (16, 17, 'sp4_h_r_33')
// (17, 13, 'sp4_r_v_b_41')
// (17, 14, 'sp4_r_v_b_28')
// (17, 14, 'sp4_r_v_b_44')
// (17, 15, 'neigh_op_tnr_2')
// (17, 15, 'sp4_r_v_b_17')
// (17, 15, 'sp4_r_v_b_33')
// (17, 16, 'neigh_op_rgt_2')
// (17, 16, 'sp12_h_r_11')
// (17, 16, 'sp4_h_r_7')
// (17, 16, 'sp4_r_v_b_20')
// (17, 16, 'sp4_r_v_b_4')
// (17, 17, 'local_g0_2')
// (17, 17, 'lutff_7/in_1')
// (17, 17, 'neigh_op_bnr_2')
// (17, 17, 'sp4_h_r_44')
// (17, 17, 'sp4_r_v_b_9')
// (18, 12, 'sp4_v_t_41')
// (18, 13, 'local_g2_1')
// (18, 13, 'lutff_4/in_1')
// (18, 13, 'sp4_v_b_41')
// (18, 13, 'sp4_v_t_44')
// (18, 14, 'local_g3_4')
// (18, 14, 'lutff_0/in_1')
// (18, 14, 'sp4_r_v_b_45')
// (18, 14, 'sp4_v_b_28')
// (18, 14, 'sp4_v_b_44')
// (18, 15, 'neigh_op_top_2')
// (18, 15, 'sp4_r_v_b_32')
// (18, 15, 'sp4_v_b_17')
// (18, 15, 'sp4_v_b_33')
// (18, 16, 'local_g1_2')
// (18, 16, 'lutff_2/in_1')
// (18, 16, 'lutff_2/out')
// (18, 16, 'sp12_h_r_12')
// (18, 16, 'sp4_h_r_18')
// (18, 16, 'sp4_r_v_b_21')
// (18, 16, 'sp4_v_b_20')
// (18, 16, 'sp4_v_b_4')
// (18, 17, 'neigh_op_bot_2')
// (18, 17, 'sp4_h_l_44')
// (18, 17, 'sp4_r_v_b_8')
// (18, 17, 'sp4_v_b_9')
// (19, 13, 'sp4_v_t_45')
// (19, 14, 'sp4_v_b_45')
// (19, 15, 'neigh_op_tnl_2')
// (19, 15, 'sp4_v_b_32')
// (19, 16, 'neigh_op_lft_2')
// (19, 16, 'sp12_h_r_15')
// (19, 16, 'sp4_h_r_31')
// (19, 16, 'sp4_v_b_21')
// (19, 17, 'local_g2_2')
// (19, 17, 'lutff_6/in_0')
// (19, 17, 'neigh_op_bnl_2')
// (19, 17, 'sp4_h_r_2')
// (19, 17, 'sp4_v_b_8')
// (20, 13, 'sp4_r_v_b_38')
// (20, 14, 'local_g1_3')
// (20, 14, 'lutff_5/in_3')
// (20, 14, 'sp4_r_v_b_27')
// (20, 15, 'sp4_r_v_b_14')
// (20, 16, 'sp12_h_r_16')
// (20, 16, 'sp4_h_r_42')
// (20, 16, 'sp4_r_v_b_3')
// (20, 17, 'sp4_h_r_15')
// (20, 17, 'sp4_r_v_b_37')
// (20, 18, 'sp4_r_v_b_24')
// (20, 19, 'sp4_r_v_b_13')
// (20, 20, 'sp4_r_v_b_0')
// (21, 12, 'sp4_v_t_38')
// (21, 13, 'sp4_v_b_38')
// (21, 14, 'sp4_v_b_27')
// (21, 15, 'sp4_v_b_14')
// (21, 16, 'sp12_h_r_19')
// (21, 16, 'sp4_h_l_42')
// (21, 16, 'sp4_h_r_10')
// (21, 16, 'sp4_v_b_3')
// (21, 16, 'sp4_v_t_37')
// (21, 17, 'sp4_h_r_26')
// (21, 17, 'sp4_v_b_37')
// (21, 18, 'sp4_v_b_24')
// (21, 19, 'local_g0_5')
// (21, 19, 'lutff_2/in_1')
// (21, 19, 'sp4_v_b_13')
// (21, 20, 'sp4_v_b_0')
// (22, 16, 'sp12_h_r_20')
// (22, 16, 'sp4_h_r_23')
// (22, 17, 'local_g2_7')
// (22, 17, 'lutff_6/in_1')
// (22, 17, 'sp4_h_r_39')
// (22, 18, 'local_g2_7')
// (22, 18, 'lutff_6/in_1')
// (22, 18, 'sp4_r_v_b_39')
// (22, 19, 'sp4_r_v_b_26')
// (22, 20, 'sp4_r_v_b_15')
// (22, 21, 'sp4_r_v_b_2')
// (23, 16, 'sp12_h_r_23')
// (23, 16, 'sp4_h_r_34')
// (23, 17, 'sp4_h_l_39')
// (23, 17, 'sp4_v_t_39')
// (23, 18, 'sp4_v_b_39')
// (23, 19, 'sp4_v_b_26')
// (23, 20, 'sp4_v_b_15')
// (23, 21, 'sp4_v_b_2')
// (24, 16, 'sp12_h_l_23')
// (24, 16, 'sp4_h_r_47')
// (25, 16, 'sp4_h_l_47')

wire n596;
// (12, 16, 'sp4_h_r_7')
// (13, 13, 'sp4_h_r_7')
// (13, 16, 'sp4_h_r_18')
// (14, 13, 'sp4_h_r_18')
// (14, 16, 'sp4_h_r_31')
// (15, 12, 'neigh_op_tnr_5')
// (15, 13, 'neigh_op_rgt_5')
// (15, 13, 'sp4_h_r_31')
// (15, 13, 'sp4_r_v_b_42')
// (15, 14, 'neigh_op_bnr_5')
// (15, 14, 'sp4_r_v_b_31')
// (15, 15, 'sp4_r_v_b_18')
// (15, 16, 'sp4_h_r_42')
// (15, 16, 'sp4_r_v_b_7')
// (16, 12, 'neigh_op_top_5')
// (16, 12, 'sp4_h_r_0')
// (16, 12, 'sp4_v_t_42')
// (16, 13, 'lutff_5/out')
// (16, 13, 'sp4_h_r_42')
// (16, 13, 'sp4_r_v_b_43')
// (16, 13, 'sp4_v_b_42')
// (16, 14, 'neigh_op_bot_5')
// (16, 14, 'sp4_r_v_b_30')
// (16, 14, 'sp4_v_b_31')
// (16, 15, 'sp4_r_v_b_19')
// (16, 15, 'sp4_v_b_18')
// (16, 16, 'sp4_h_l_42')
// (16, 16, 'sp4_h_r_10')
// (16, 16, 'sp4_h_r_3')
// (16, 16, 'sp4_r_v_b_6')
// (16, 16, 'sp4_v_b_7')
// (17, 12, 'neigh_op_tnl_5')
// (17, 12, 'sp4_h_r_13')
// (17, 12, 'sp4_h_r_6')
// (17, 12, 'sp4_v_t_43')
// (17, 13, 'local_g0_2')
// (17, 13, 'lutff_global/cen')
// (17, 13, 'neigh_op_lft_5')
// (17, 13, 'sp4_h_l_42')
// (17, 13, 'sp4_h_r_10')
// (17, 13, 'sp4_v_b_43')
// (17, 14, 'neigh_op_bnl_5')
// (17, 14, 'sp4_v_b_30')
// (17, 15, 'sp4_v_b_19')
// (17, 16, 'sp4_h_r_14')
// (17, 16, 'sp4_h_r_23')
// (17, 16, 'sp4_v_b_6')
// (18, 12, 'sp4_h_r_19')
// (18, 12, 'sp4_h_r_24')
// (18, 13, 'sp4_h_r_23')
// (18, 16, 'sp4_h_r_27')
// (18, 16, 'sp4_h_r_34')
// (19, 9, 'local_g3_3')
// (19, 9, 'lutff_global/cen')
// (19, 9, 'sp4_r_v_b_43')
// (19, 10, 'sp4_r_v_b_30')
// (19, 11, 'sp4_r_v_b_19')
// (19, 12, 'sp4_h_r_30')
// (19, 12, 'sp4_h_r_37')
// (19, 12, 'sp4_r_v_b_6')
// (19, 13, 'local_g2_2')
// (19, 13, 'lutff_global/cen')
// (19, 13, 'sp4_h_r_34')
// (19, 13, 'sp4_r_v_b_44')
// (19, 14, 'local_g0_2')
// (19, 14, 'lutff_global/cen')
// (19, 14, 'sp4_r_v_b_33')
// (19, 15, 'sp4_r_v_b_20')
// (19, 16, 'sp4_h_r_38')
// (19, 16, 'sp4_h_r_47')
// (19, 16, 'sp4_r_v_b_9')
// (19, 17, 'sp4_r_v_b_47')
// (19, 18, 'local_g2_2')
// (19, 18, 'lutff_global/cen')
// (19, 18, 'sp4_r_v_b_34')
// (19, 19, 'sp4_r_v_b_23')
// (19, 20, 'sp4_r_v_b_10')
// (20, 8, 'sp4_v_t_43')
// (20, 9, 'sp4_v_b_43')
// (20, 10, 'sp4_v_b_30')
// (20, 11, 'sp4_v_b_19')
// (20, 12, 'sp4_h_l_37')
// (20, 12, 'sp4_h_r_43')
// (20, 12, 'sp4_v_b_6')
// (20, 12, 'sp4_v_t_44')
// (20, 13, 'sp4_h_r_47')
// (20, 13, 'sp4_r_v_b_43')
// (20, 13, 'sp4_v_b_44')
// (20, 14, 'sp4_r_v_b_30')
// (20, 14, 'sp4_v_b_33')
// (20, 15, 'sp4_r_v_b_19')
// (20, 15, 'sp4_v_b_20')
// (20, 16, 'sp4_h_l_38')
// (20, 16, 'sp4_h_l_47')
// (20, 16, 'sp4_h_r_10')
// (20, 16, 'sp4_h_r_6')
// (20, 16, 'sp4_r_v_b_6')
// (20, 16, 'sp4_v_b_9')
// (20, 16, 'sp4_v_t_47')
// (20, 17, 'sp4_v_b_47')
// (20, 18, 'sp4_v_b_34')
// (20, 19, 'sp4_v_b_23')
// (20, 20, 'sp4_v_b_10')
// (21, 12, 'sp4_h_l_43')
// (21, 12, 'sp4_v_t_43')
// (21, 13, 'local_g3_3')
// (21, 13, 'lutff_global/cen')
// (21, 13, 'sp4_h_l_47')
// (21, 13, 'sp4_v_b_43')
// (21, 14, 'sp4_v_b_30')
// (21, 15, 'sp4_v_b_19')
// (21, 16, 'local_g1_3')
// (21, 16, 'lutff_global/cen')
// (21, 16, 'sp4_h_r_19')
// (21, 16, 'sp4_h_r_23')
// (21, 16, 'sp4_v_b_6')
// (22, 16, 'local_g2_2')
// (22, 16, 'lutff_global/cen')
// (22, 16, 'sp4_h_r_30')
// (22, 16, 'sp4_h_r_34')
// (23, 16, 'sp4_h_r_43')
// (23, 16, 'sp4_h_r_47')
// (24, 16, 'sp4_h_l_43')
// (24, 16, 'sp4_h_l_47')

wire n597;
// (12, 17, 'lutff_0/cout')
// (12, 17, 'lutff_1/in_3')

wire n598;
// (12, 17, 'lutff_1/cout')
// (12, 17, 'lutff_2/in_3')

wire n599;
// (12, 17, 'lutff_2/cout')
// (12, 17, 'lutff_3/in_3')

wire n600;
// (12, 17, 'lutff_3/cout')
// (12, 17, 'lutff_4/in_3')

wire n601;
// (12, 17, 'lutff_4/cout')
// (12, 17, 'lutff_5/in_3')

wire n602;
// (12, 17, 'lutff_5/cout')
// (12, 17, 'lutff_6/in_3')

wire n603;
// (12, 17, 'lutff_6/cout')
// (12, 17, 'lutff_7/in_3')

wire n604;
// (12, 17, 'lutff_7/cout')
// (12, 18, 'carry_in')
// (12, 18, 'carry_in_mux')
// (12, 18, 'lutff_0/in_3')

wire n605;
// (12, 17, 'neigh_op_tnr_4')
// (12, 18, 'neigh_op_rgt_4')
// (12, 19, 'neigh_op_bnr_4')
// (13, 17, 'neigh_op_top_4')
// (13, 18, 'local_g0_4')
// (13, 18, 'lutff_4/in_2')
// (13, 18, 'lutff_4/out')
// (13, 18, 'sp12_h_r_0')
// (13, 19, 'neigh_op_bot_4')
// (14, 17, 'neigh_op_tnl_4')
// (14, 18, 'neigh_op_lft_4')
// (14, 18, 'sp12_h_r_3')
// (14, 19, 'neigh_op_bnl_4')
// (15, 18, 'sp12_h_r_4')
// (16, 18, 'sp12_h_r_7')
// (17, 18, 'local_g0_0')
// (17, 18, 'lutff_4/in_2')
// (17, 18, 'sp12_h_r_8')
// (18, 18, 'sp12_h_r_11')
// (19, 18, 'sp12_h_r_12')
// (20, 18, 'sp12_h_r_15')
// (21, 18, 'sp12_h_r_16')
// (22, 18, 'sp12_h_r_19')
// (23, 18, 'sp12_h_r_20')
// (24, 18, 'sp12_h_r_23')
// (25, 18, 'sp12_h_l_23')

wire n606;
// (12, 17, 'neigh_op_tnr_5')
// (12, 18, 'neigh_op_rgt_5')
// (12, 18, 'sp12_h_r_1')
// (12, 19, 'neigh_op_bnr_5')
// (13, 17, 'neigh_op_top_5')
// (13, 18, 'local_g1_2')
// (13, 18, 'lutff_5/in_2')
// (13, 18, 'lutff_5/out')
// (13, 18, 'sp12_h_r_2')
// (13, 19, 'neigh_op_bot_5')
// (14, 17, 'neigh_op_tnl_5')
// (14, 18, 'neigh_op_lft_5')
// (14, 18, 'sp12_h_r_5')
// (14, 19, 'neigh_op_bnl_5')
// (15, 18, 'sp12_h_r_6')
// (16, 18, 'sp12_h_r_9')
// (17, 18, 'local_g1_2')
// (17, 18, 'lutff_5/in_2')
// (17, 18, 'sp12_h_r_10')
// (18, 18, 'sp12_h_r_13')
// (19, 18, 'sp12_h_r_14')
// (20, 18, 'sp12_h_r_17')
// (21, 18, 'sp12_h_r_18')
// (22, 18, 'sp12_h_r_21')
// (23, 18, 'sp12_h_r_22')
// (24, 18, 'sp12_h_l_22')

wire n607;
// (12, 17, 'sp12_h_r_0')
// (13, 17, 'sp12_h_r_3')
// (14, 17, 'local_g0_4')
// (14, 17, 'lutff_3/in_3')
// (14, 17, 'sp12_h_r_4')
// (15, 17, 'sp12_h_r_7')
// (16, 17, 'sp12_h_r_8')
// (17, 16, 'neigh_op_tnr_2')
// (17, 17, 'neigh_op_rgt_2')
// (17, 17, 'sp12_h_r_11')
// (17, 18, 'neigh_op_bnr_2')
// (18, 16, 'neigh_op_top_2')
// (18, 17, 'lutff_2/out')
// (18, 17, 'sp12_h_r_12')
// (18, 18, 'neigh_op_bot_2')
// (19, 16, 'neigh_op_tnl_2')
// (19, 17, 'neigh_op_lft_2')
// (19, 17, 'sp12_h_r_15')
// (19, 18, 'neigh_op_bnl_2')
// (20, 17, 'sp12_h_r_16')
// (21, 17, 'sp12_h_r_19')
// (22, 17, 'sp12_h_r_20')
// (23, 17, 'sp12_h_r_23')
// (24, 17, 'sp12_h_l_23')

wire n608;
// (12, 17, 'sp12_h_r_1')
// (13, 17, 'sp12_h_r_2')
// (14, 17, 'sp12_h_r_5')
// (15, 17, 'sp12_h_r_6')
// (16, 17, 'sp12_h_r_9')
// (17, 17, 'sp12_h_r_10')
// (18, 17, 'sp12_h_r_13')
// (19, 17, 'local_g0_6')
// (19, 17, 'lutff_3/in_3')
// (19, 17, 'sp12_h_r_14')
// (20, 17, 'sp12_h_r_17')
// (21, 17, 'sp12_h_r_18')
// (22, 16, 'neigh_op_tnr_7')
// (22, 17, 'neigh_op_rgt_7')
// (22, 17, 'sp12_h_r_21')
// (22, 18, 'neigh_op_bnr_7')
// (23, 16, 'neigh_op_top_7')
// (23, 17, 'lutff_7/out')
// (23, 17, 'sp12_h_r_22')
// (23, 18, 'neigh_op_bot_7')
// (24, 16, 'neigh_op_tnl_7')
// (24, 17, 'neigh_op_lft_7')
// (24, 17, 'sp12_h_l_22')
// (24, 18, 'neigh_op_bnl_7')

wire n609;
// (12, 17, 'sp4_h_r_7')
// (13, 17, 'sp4_h_r_18')
// (14, 17, 'sp4_h_r_31')
// (15, 13, 'neigh_op_tnr_4')
// (15, 14, 'neigh_op_rgt_4')
// (15, 14, 'sp4_r_v_b_40')
// (15, 15, 'neigh_op_bnr_4')
// (15, 15, 'sp4_r_v_b_29')
// (15, 16, 'sp4_r_v_b_16')
// (15, 17, 'local_g2_2')
// (15, 17, 'lutff_global/cen')
// (15, 17, 'sp4_h_r_42')
// (15, 17, 'sp4_r_v_b_5')
// (16, 13, 'neigh_op_top_4')
// (16, 13, 'sp4_v_t_40')
// (16, 14, 'lutff_4/out')
// (16, 14, 'sp4_v_b_40')
// (16, 15, 'neigh_op_bot_4')
// (16, 15, 'sp4_v_b_29')
// (16, 16, 'sp4_v_b_16')
// (16, 17, 'sp4_h_l_42')
// (16, 17, 'sp4_h_r_11')
// (16, 17, 'sp4_v_b_5')
// (17, 13, 'neigh_op_tnl_4')
// (17, 14, 'neigh_op_lft_4')
// (17, 15, 'neigh_op_bnl_4')
// (17, 17, 'sp4_h_r_22')
// (18, 17, 'sp4_h_r_35')
// (19, 17, 'sp4_h_r_46')
// (20, 17, 'sp4_h_l_46')

wire n610;
// (12, 18, 'lutff_0/cout')
// (12, 18, 'lutff_1/in_3')

wire n611;
// (12, 18, 'lutff_1/cout')
// (12, 18, 'lutff_2/in_3')

wire n612;
// (12, 18, 'lutff_2/cout')
// (12, 18, 'lutff_3/in_3')

wire n613;
// (12, 18, 'lutff_3/cout')
// (12, 18, 'lutff_4/in_3')

wire n614;
// (12, 18, 'lutff_4/cout')
// (12, 18, 'lutff_5/in_3')

wire n615;
// (12, 18, 'lutff_5/cout')
// (12, 18, 'lutff_6/in_3')

wire n616;
// (12, 18, 'lutff_6/cout')
// (12, 18, 'lutff_7/in_3')

wire n617;
// (12, 18, 'neigh_op_tnr_4')
// (12, 19, 'neigh_op_rgt_4')
// (12, 20, 'neigh_op_bnr_4')
// (13, 18, 'neigh_op_top_4')
// (13, 19, 'local_g0_4')
// (13, 19, 'lutff_4/in_2')
// (13, 19, 'lutff_4/out')
// (13, 19, 'sp12_h_r_0')
// (13, 20, 'neigh_op_bot_4')
// (14, 18, 'neigh_op_tnl_4')
// (14, 19, 'neigh_op_lft_4')
// (14, 19, 'sp12_h_r_3')
// (14, 20, 'neigh_op_bnl_4')
// (15, 19, 'sp12_h_r_4')
// (16, 19, 'sp12_h_r_7')
// (17, 19, 'local_g0_0')
// (17, 19, 'lutff_4/in_2')
// (17, 19, 'sp12_h_r_8')
// (18, 19, 'sp12_h_r_11')
// (19, 19, 'sp12_h_r_12')
// (20, 19, 'sp12_h_r_15')
// (21, 19, 'sp12_h_r_16')
// (22, 19, 'sp12_h_r_19')
// (23, 19, 'sp12_h_r_20')
// (24, 19, 'sp12_h_r_23')
// (25, 19, 'sp12_h_l_23')

wire n618;
// (12, 18, 'neigh_op_tnr_5')
// (12, 19, 'neigh_op_rgt_5')
// (12, 19, 'sp12_h_r_1')
// (12, 20, 'neigh_op_bnr_5')
// (13, 18, 'neigh_op_top_5')
// (13, 19, 'local_g0_2')
// (13, 19, 'lutff_5/in_1')
// (13, 19, 'lutff_5/out')
// (13, 19, 'sp12_h_r_2')
// (13, 20, 'neigh_op_bot_5')
// (14, 18, 'neigh_op_tnl_5')
// (14, 19, 'neigh_op_lft_5')
// (14, 19, 'sp12_h_r_5')
// (14, 20, 'neigh_op_bnl_5')
// (15, 19, 'sp12_h_r_6')
// (16, 19, 'sp12_h_r_9')
// (17, 19, 'local_g1_2')
// (17, 19, 'lutff_5/in_2')
// (17, 19, 'sp12_h_r_10')
// (18, 19, 'sp12_h_r_13')
// (19, 19, 'sp12_h_r_14')
// (20, 19, 'sp12_h_r_17')
// (21, 19, 'sp12_h_r_18')
// (22, 19, 'sp12_h_r_21')
// (23, 19, 'sp12_h_r_22')
// (24, 19, 'sp12_h_l_22')

wire n619;
// (12, 18, 'sp4_h_r_10')
// (13, 18, 'sp4_h_r_23')
// (14, 13, 'sp4_r_v_b_47')
// (14, 14, 'sp4_r_v_b_34')
// (14, 15, 'sp4_r_v_b_23')
// (14, 16, 'sp4_r_v_b_10')
// (14, 17, 'sp4_r_v_b_42')
// (14, 18, 'sp4_h_r_34')
// (14, 18, 'sp4_r_v_b_31')
// (14, 19, 'sp4_r_v_b_18')
// (14, 20, 'sp4_r_v_b_7')
// (15, 12, 'sp4_h_r_10')
// (15, 12, 'sp4_v_t_47')
// (15, 13, 'sp4_v_b_47')
// (15, 14, 'sp4_v_b_34')
// (15, 15, 'sp4_v_b_23')
// (15, 16, 'sp4_v_b_10')
// (15, 16, 'sp4_v_t_42')
// (15, 17, 'sp4_v_b_42')
// (15, 18, 'sp4_h_r_47')
// (15, 18, 'sp4_r_v_b_42')
// (15, 18, 'sp4_v_b_31')
// (15, 19, 'neigh_op_tnr_1')
// (15, 19, 'sp4_r_v_b_31')
// (15, 19, 'sp4_r_v_b_47')
// (15, 19, 'sp4_v_b_18')
// (15, 20, 'neigh_op_rgt_1')
// (15, 20, 'sp4_h_r_7')
// (15, 20, 'sp4_r_v_b_18')
// (15, 20, 'sp4_r_v_b_34')
// (15, 20, 'sp4_v_b_7')
// (15, 21, 'neigh_op_bnr_1')
// (15, 21, 'sp4_r_v_b_23')
// (15, 21, 'sp4_r_v_b_7')
// (15, 22, 'sp4_r_v_b_10')
// (16, 12, 'sp4_h_r_23')
// (16, 17, 'sp4_h_r_7')
// (16, 17, 'sp4_v_t_42')
// (16, 18, 'sp4_h_l_47')
// (16, 18, 'sp4_h_r_6')
// (16, 18, 'sp4_v_b_42')
// (16, 18, 'sp4_v_t_47')
// (16, 19, 'neigh_op_top_1')
// (16, 19, 'sp4_v_b_31')
// (16, 19, 'sp4_v_b_47')
// (16, 20, 'lutff_1/out')
// (16, 20, 'sp4_h_r_18')
// (16, 20, 'sp4_v_b_18')
// (16, 20, 'sp4_v_b_34')
// (16, 21, 'neigh_op_bot_1')
// (16, 21, 'sp4_v_b_23')
// (16, 21, 'sp4_v_b_7')
// (16, 22, 'sp4_v_b_10')
// (17, 12, 'local_g2_2')
// (17, 12, 'lutff_global/cen')
// (17, 12, 'sp4_h_r_34')
// (17, 17, 'sp4_h_r_18')
// (17, 18, 'sp4_h_r_19')
// (17, 19, 'neigh_op_tnl_1')
// (17, 20, 'neigh_op_lft_1')
// (17, 20, 'sp4_h_r_31')
// (17, 21, 'neigh_op_bnl_1')
// (18, 12, 'sp4_h_r_47')
// (18, 17, 'sp4_h_r_31')
// (18, 18, 'sp4_h_r_30')
// (18, 20, 'sp4_h_r_42')
// (19, 12, 'sp4_h_l_47')
// (19, 15, 'local_g3_3')
// (19, 15, 'lutff_global/cen')
// (19, 15, 'sp4_r_v_b_43')
// (19, 16, 'sp4_r_v_b_30')
// (19, 17, 'sp4_h_r_42')
// (19, 17, 'sp4_r_v_b_19')
// (19, 18, 'sp4_h_r_43')
// (19, 18, 'sp4_r_v_b_6')
// (19, 20, 'sp4_h_l_42')
// (20, 14, 'sp4_v_t_43')
// (20, 15, 'sp4_v_b_43')
// (20, 16, 'sp4_v_b_30')
// (20, 17, 'sp4_h_l_42')
// (20, 17, 'sp4_h_r_7')
// (20, 17, 'sp4_v_b_19')
// (20, 18, 'sp4_h_l_43')
// (20, 18, 'sp4_h_r_2')
// (20, 18, 'sp4_v_b_6')
// (21, 17, 'sp4_h_r_18')
// (21, 18, 'sp4_h_r_15')
// (22, 17, 'sp4_h_r_31')
// (22, 18, 'sp4_h_r_26')
// (23, 15, 'sp4_r_v_b_39')
// (23, 16, 'sp4_r_v_b_26')
// (23, 17, 'local_g2_2')
// (23, 17, 'lutff_global/cen')
// (23, 17, 'sp4_h_r_42')
// (23, 17, 'sp4_r_v_b_15')
// (23, 18, 'sp4_h_r_39')
// (23, 18, 'sp4_r_v_b_2')
// (24, 14, 'sp4_v_t_39')
// (24, 15, 'sp4_v_b_39')
// (24, 16, 'local_g2_2')
// (24, 16, 'lutff_global/cen')
// (24, 16, 'sp4_v_b_26')
// (24, 17, 'sp4_h_l_42')
// (24, 17, 'sp4_v_b_15')
// (24, 18, 'sp4_h_l_39')
// (24, 18, 'sp4_v_b_2')

wire n620;
// (12, 19, 'local_g0_2')
// (12, 19, 'lutff_global/cen')
// (12, 19, 'sp4_h_r_2')
// (13, 19, 'sp4_h_r_15')
// (14, 15, 'neigh_op_tnr_3')
// (14, 16, 'neigh_op_rgt_3')
// (14, 17, 'neigh_op_bnr_3')
// (14, 19, 'sp4_h_r_26')
// (15, 15, 'neigh_op_top_3')
// (15, 16, 'lutff_3/out')
// (15, 16, 'sp4_r_v_b_39')
// (15, 17, 'neigh_op_bot_3')
// (15, 17, 'sp4_r_v_b_26')
// (15, 18, 'sp4_r_v_b_15')
// (15, 19, 'sp4_h_r_39')
// (15, 19, 'sp4_r_v_b_2')
// (16, 15, 'neigh_op_tnl_3')
// (16, 15, 'sp4_v_t_39')
// (16, 16, 'neigh_op_lft_3')
// (16, 16, 'sp4_v_b_39')
// (16, 17, 'neigh_op_bnl_3')
// (16, 17, 'sp4_v_b_26')
// (16, 18, 'sp4_v_b_15')
// (16, 19, 'sp4_h_l_39')
// (16, 19, 'sp4_v_b_2')

wire n621;
// (12, 19, 'neigh_op_tnr_0')
// (12, 20, 'neigh_op_rgt_0')
// (12, 21, 'neigh_op_bnr_0')
// (13, 19, 'neigh_op_top_0')
// (13, 20, 'local_g1_0')
// (13, 20, 'lutff_0/in_1')
// (13, 20, 'lutff_0/out')
// (13, 21, 'neigh_op_bot_0')
// (14, 19, 'neigh_op_tnl_0')
// (14, 20, 'neigh_op_lft_0')
// (14, 21, 'neigh_op_bnl_0')

wire n622;
// (12, 19, 'neigh_op_tnr_1')
// (12, 20, 'neigh_op_rgt_1')
// (12, 21, 'neigh_op_bnr_1')
// (13, 19, 'neigh_op_top_1')
// (13, 20, 'local_g3_1')
// (13, 20, 'lutff_1/in_1')
// (13, 20, 'lutff_1/out')
// (13, 21, 'neigh_op_bot_1')
// (14, 19, 'neigh_op_tnl_1')
// (14, 20, 'neigh_op_lft_1')
// (14, 21, 'neigh_op_bnl_1')

wire n623;
// (12, 19, 'neigh_op_tnr_2')
// (12, 20, 'neigh_op_rgt_2')
// (12, 21, 'neigh_op_bnr_2')
// (13, 19, 'neigh_op_top_2')
// (13, 20, 'local_g1_2')
// (13, 20, 'lutff_2/in_1')
// (13, 20, 'lutff_2/out')
// (13, 21, 'neigh_op_bot_2')
// (14, 19, 'neigh_op_tnl_2')
// (14, 20, 'neigh_op_lft_2')
// (14, 21, 'neigh_op_bnl_2')

wire n624;
// (12, 19, 'neigh_op_tnr_3')
// (12, 20, 'neigh_op_rgt_3')
// (12, 21, 'neigh_op_bnr_3')
// (13, 19, 'neigh_op_top_3')
// (13, 20, 'local_g1_3')
// (13, 20, 'lutff_3/in_1')
// (13, 20, 'lutff_3/out')
// (13, 21, 'neigh_op_bot_3')
// (14, 19, 'neigh_op_tnl_3')
// (14, 20, 'neigh_op_lft_3')
// (14, 21, 'neigh_op_bnl_3')

wire n625;
// (12, 19, 'neigh_op_tnr_4')
// (12, 20, 'neigh_op_rgt_4')
// (12, 21, 'neigh_op_bnr_4')
// (13, 19, 'neigh_op_top_4')
// (13, 20, 'local_g1_4')
// (13, 20, 'lutff_4/in_1')
// (13, 20, 'lutff_4/out')
// (13, 21, 'neigh_op_bot_4')
// (14, 19, 'neigh_op_tnl_4')
// (14, 20, 'neigh_op_lft_4')
// (14, 21, 'neigh_op_bnl_4')

wire n626;
// (12, 19, 'neigh_op_tnr_5')
// (12, 20, 'neigh_op_rgt_5')
// (12, 21, 'neigh_op_bnr_5')
// (13, 19, 'neigh_op_top_5')
// (13, 20, 'local_g1_5')
// (13, 20, 'lutff_5/in_1')
// (13, 20, 'lutff_5/out')
// (13, 21, 'neigh_op_bot_5')
// (14, 19, 'neigh_op_tnl_5')
// (14, 20, 'neigh_op_lft_5')
// (14, 21, 'neigh_op_bnl_5')

wire n627;
// (12, 19, 'neigh_op_tnr_6')
// (12, 20, 'neigh_op_rgt_6')
// (12, 21, 'neigh_op_bnr_6')
// (13, 19, 'neigh_op_top_6')
// (13, 20, 'local_g1_6')
// (13, 20, 'lutff_6/in_1')
// (13, 20, 'lutff_6/out')
// (13, 21, 'neigh_op_bot_6')
// (14, 19, 'neigh_op_tnl_6')
// (14, 20, 'neigh_op_lft_6')
// (14, 21, 'neigh_op_bnl_6')

wire n628;
// (12, 19, 'neigh_op_tnr_7')
// (12, 20, 'neigh_op_rgt_7')
// (12, 21, 'neigh_op_bnr_7')
// (13, 19, 'neigh_op_top_7')
// (13, 20, 'local_g3_7')
// (13, 20, 'lutff_7/in_1')
// (13, 20, 'lutff_7/out')
// (13, 21, 'neigh_op_bot_7')
// (14, 19, 'neigh_op_tnl_7')
// (14, 20, 'neigh_op_lft_7')
// (14, 21, 'neigh_op_bnl_7')

wire n629;
// (12, 19, 'sp4_h_r_7')
// (13, 19, 'sp4_h_r_18')
// (14, 19, 'sp4_h_r_31')
// (14, 21, 'local_g3_3')
// (14, 21, 'lutff_global/cen')
// (14, 21, 'sp4_r_v_b_43')
// (14, 22, 'sp4_r_v_b_30')
// (14, 23, 'sp4_r_v_b_19')
// (14, 24, 'sp4_r_v_b_6')
// (15, 19, 'local_g2_2')
// (15, 19, 'lutff_global/cen')
// (15, 19, 'neigh_op_tnr_5')
// (15, 19, 'sp4_h_r_42')
// (15, 20, 'neigh_op_rgt_5')
// (15, 20, 'sp12_h_r_1')
// (15, 20, 'sp4_h_r_0')
// (15, 20, 'sp4_r_v_b_42')
// (15, 20, 'sp4_v_t_43')
// (15, 21, 'neigh_op_bnr_5')
// (15, 21, 'sp4_r_v_b_31')
// (15, 21, 'sp4_v_b_43')
// (15, 22, 'sp4_r_v_b_18')
// (15, 22, 'sp4_v_b_30')
// (15, 23, 'sp4_r_v_b_7')
// (15, 23, 'sp4_v_b_19')
// (15, 24, 'sp4_v_b_6')
// (16, 19, 'neigh_op_top_5')
// (16, 19, 'sp4_h_l_42')
// (16, 19, 'sp4_v_t_42')
// (16, 20, 'lutff_5/out')
// (16, 20, 'sp12_h_r_2')
// (16, 20, 'sp4_h_r_13')
// (16, 20, 'sp4_v_b_42')
// (16, 21, 'neigh_op_bot_5')
// (16, 21, 'sp4_v_b_31')
// (16, 22, 'sp4_v_b_18')
// (16, 23, 'sp4_v_b_7')
// (17, 19, 'neigh_op_tnl_5')
// (17, 20, 'neigh_op_lft_5')
// (17, 20, 'sp12_h_r_5')
// (17, 20, 'sp4_h_r_24')
// (17, 21, 'neigh_op_bnl_5')
// (18, 20, 'sp12_h_r_6')
// (18, 20, 'sp4_h_r_37')
// (19, 20, 'sp12_h_r_9')
// (19, 20, 'sp4_h_l_37')
// (20, 20, 'sp12_h_r_10')
// (21, 20, 'sp12_h_r_13')
// (22, 20, 'sp12_h_r_14')
// (23, 20, 'sp12_h_r_17')
// (24, 20, 'sp12_h_r_18')
// (25, 20, 'sp12_h_r_21')
// (26, 20, 'sp12_h_r_22')
// (27, 20, 'sp12_h_l_22')

wire n630;
// (12, 19, 'sp4_r_v_b_38')
// (12, 20, 'neigh_op_tnr_7')
// (12, 20, 'sp4_r_v_b_27')
// (12, 21, 'neigh_op_rgt_7')
// (12, 21, 'sp4_r_v_b_14')
// (12, 22, 'neigh_op_bnr_7')
// (12, 22, 'sp4_r_v_b_3')
// (13, 18, 'sp4_h_r_8')
// (13, 18, 'sp4_v_t_38')
// (13, 19, 'sp4_r_v_b_39')
// (13, 19, 'sp4_v_b_38')
// (13, 20, 'neigh_op_top_7')
// (13, 20, 'sp4_r_v_b_26')
// (13, 20, 'sp4_v_b_27')
// (13, 21, 'lutff_7/out')
// (13, 21, 'sp4_r_v_b_15')
// (13, 21, 'sp4_v_b_14')
// (13, 22, 'neigh_op_bot_7')
// (13, 22, 'sp4_r_v_b_2')
// (13, 22, 'sp4_v_b_3')
// (14, 18, 'local_g0_5')
// (14, 18, 'local_g1_7')
// (14, 18, 'lutff_0/in_0')
// (14, 18, 'lutff_1/in_0')
// (14, 18, 'lutff_2/in_0')
// (14, 18, 'lutff_3/in_0')
// (14, 18, 'lutff_4/in_0')
// (14, 18, 'lutff_5/in_0')
// (14, 18, 'lutff_6/in_0')
// (14, 18, 'lutff_7/in_0')
// (14, 18, 'sp4_h_r_21')
// (14, 18, 'sp4_h_r_7')
// (14, 18, 'sp4_v_t_39')
// (14, 19, 'local_g2_7')
// (14, 19, 'local_g3_7')
// (14, 19, 'lutff_0/in_0')
// (14, 19, 'lutff_1/in_0')
// (14, 19, 'lutff_2/in_0')
// (14, 19, 'lutff_3/in_0')
// (14, 19, 'lutff_4/in_0')
// (14, 19, 'lutff_5/in_0')
// (14, 19, 'lutff_6/in_0')
// (14, 19, 'lutff_7/in_0')
// (14, 19, 'sp4_v_b_39')
// (14, 20, 'local_g2_7')
// (14, 20, 'local_g3_7')
// (14, 20, 'lutff_0/in_0')
// (14, 20, 'lutff_1/in_0')
// (14, 20, 'lutff_2/in_0')
// (14, 20, 'lutff_3/in_0')
// (14, 20, 'lutff_4/in_0')
// (14, 20, 'lutff_5/in_0')
// (14, 20, 'lutff_6/in_0')
// (14, 20, 'lutff_7/in_0')
// (14, 20, 'neigh_op_tnl_7')
// (14, 20, 'sp4_v_b_26')
// (14, 21, 'neigh_op_lft_7')
// (14, 21, 'sp4_v_b_15')
// (14, 22, 'neigh_op_bnl_7')
// (14, 22, 'sp4_v_b_2')
// (15, 18, 'sp4_h_r_18')
// (15, 18, 'sp4_h_r_32')
// (16, 18, 'sp4_h_r_31')
// (16, 18, 'sp4_h_r_45')
// (17, 18, 'sp4_h_l_45')
// (17, 18, 'sp4_h_r_42')
// (18, 18, 'sp4_h_l_42')

wire n631;
// (12, 21, 'lutff_7/cout')
// (12, 22, 'carry_in')
// (12, 22, 'carry_in_mux')

wire n632;
// (12, 21, 'neigh_op_tnr_0')
// (12, 22, 'neigh_op_rgt_0')
// (12, 23, 'neigh_op_bnr_0')
// (13, 21, 'neigh_op_top_0')
// (13, 22, 'local_g0_0')
// (13, 22, 'lutff_0/in_2')
// (13, 22, 'lutff_0/out')
// (13, 23, 'neigh_op_bot_0')
// (14, 21, 'neigh_op_tnl_0')
// (14, 22, 'neigh_op_lft_0')
// (14, 23, 'neigh_op_bnl_0')

wire n633;
// (12, 21, 'neigh_op_tnr_1')
// (12, 22, 'neigh_op_rgt_1')
// (12, 23, 'neigh_op_bnr_1')
// (13, 21, 'neigh_op_top_1')
// (13, 22, 'local_g3_1')
// (13, 22, 'lutff_1/in_1')
// (13, 22, 'lutff_1/out')
// (13, 23, 'neigh_op_bot_1')
// (14, 21, 'neigh_op_tnl_1')
// (14, 22, 'neigh_op_lft_1')
// (14, 23, 'neigh_op_bnl_1')

wire n634;
// (12, 21, 'neigh_op_tnr_2')
// (12, 22, 'neigh_op_rgt_2')
// (12, 23, 'neigh_op_bnr_2')
// (13, 21, 'neigh_op_top_2')
// (13, 22, 'local_g1_2')
// (13, 22, 'lutff_2/in_1')
// (13, 22, 'lutff_2/out')
// (13, 23, 'neigh_op_bot_2')
// (14, 21, 'neigh_op_tnl_2')
// (14, 22, 'neigh_op_lft_2')
// (14, 23, 'neigh_op_bnl_2')

wire n635;
// (12, 21, 'neigh_op_tnr_3')
// (12, 22, 'neigh_op_rgt_3')
// (12, 23, 'neigh_op_bnr_3')
// (13, 21, 'neigh_op_top_3')
// (13, 22, 'local_g3_3')
// (13, 22, 'lutff_3/in_1')
// (13, 22, 'lutff_3/out')
// (13, 23, 'neigh_op_bot_3')
// (14, 21, 'neigh_op_tnl_3')
// (14, 22, 'neigh_op_lft_3')
// (14, 23, 'neigh_op_bnl_3')

wire n636;
// (12, 21, 'neigh_op_tnr_4')
// (12, 22, 'neigh_op_rgt_4')
// (12, 23, 'neigh_op_bnr_4')
// (13, 21, 'neigh_op_top_4')
// (13, 22, 'local_g2_4')
// (13, 22, 'lutff_4/in_2')
// (13, 22, 'lutff_4/out')
// (13, 23, 'neigh_op_bot_4')
// (14, 21, 'neigh_op_tnl_4')
// (14, 22, 'neigh_op_lft_4')
// (14, 23, 'neigh_op_bnl_4')

wire n637;
// (12, 21, 'neigh_op_tnr_5')
// (12, 22, 'neigh_op_rgt_5')
// (12, 23, 'neigh_op_bnr_5')
// (13, 21, 'neigh_op_top_5')
// (13, 22, 'local_g3_5')
// (13, 22, 'lutff_5/in_1')
// (13, 22, 'lutff_5/out')
// (13, 23, 'neigh_op_bot_5')
// (14, 21, 'neigh_op_tnl_5')
// (14, 22, 'neigh_op_lft_5')
// (14, 23, 'neigh_op_bnl_5')

wire n638;
// (12, 21, 'neigh_op_tnr_6')
// (12, 22, 'neigh_op_rgt_6')
// (12, 23, 'neigh_op_bnr_6')
// (13, 21, 'neigh_op_top_6')
// (13, 22, 'local_g1_6')
// (13, 22, 'lutff_6/in_1')
// (13, 22, 'lutff_6/out')
// (13, 23, 'neigh_op_bot_6')
// (14, 21, 'neigh_op_tnl_6')
// (14, 22, 'neigh_op_lft_6')
// (14, 23, 'neigh_op_bnl_6')

wire n639;
// (12, 21, 'neigh_op_tnr_7')
// (12, 22, 'neigh_op_rgt_7')
// (12, 23, 'neigh_op_bnr_7')
// (13, 21, 'neigh_op_top_7')
// (13, 22, 'local_g3_7')
// (13, 22, 'lutff_7/in_1')
// (13, 22, 'lutff_7/out')
// (13, 23, 'neigh_op_bot_7')
// (14, 21, 'neigh_op_tnl_7')
// (14, 22, 'neigh_op_lft_7')
// (14, 23, 'neigh_op_bnl_7')

wire n640;
// (12, 22, 'lutff_7/cout')
// (12, 23, 'carry_in')
// (12, 23, 'carry_in_mux')

wire n641;
// (12, 22, 'sp12_h_r_0')
// (13, 22, 'sp12_h_r_3')
// (14, 22, 'sp12_h_r_4')
// (15, 22, 'sp12_h_r_7')
// (16, 22, 'sp12_h_r_8')
// (17, 22, 'sp12_h_r_11')
// (18, 22, 'local_g1_4')
// (18, 22, 'lutff_4/in_1')
// (18, 22, 'sp12_h_r_12')
// (19, 21, 'local_g2_4')
// (19, 21, 'local_g3_4')
// (19, 21, 'lutff_0/in_1')
// (19, 21, 'lutff_1/in_3')
// (19, 21, 'lutff_2/in_1')
// (19, 21, 'lutff_3/in_3')
// (19, 21, 'lutff_4/in_1')
// (19, 21, 'lutff_5/in_3')
// (19, 21, 'lutff_6/in_2')
// (19, 21, 'lutff_7/in_3')
// (19, 21, 'neigh_op_tnr_4')
// (19, 22, 'neigh_op_rgt_4')
// (19, 22, 'sp12_h_r_15')
// (19, 23, 'neigh_op_bnr_4')
// (20, 21, 'neigh_op_top_4')
// (20, 22, 'local_g1_4')
// (20, 22, 'lutff_2/in_1')
// (20, 22, 'lutff_4/out')
// (20, 22, 'sp12_h_r_16')
// (20, 23, 'neigh_op_bot_4')
// (21, 21, 'neigh_op_tnl_4')
// (21, 22, 'neigh_op_lft_4')
// (21, 22, 'sp12_h_r_19')
// (21, 23, 'neigh_op_bnl_4')
// (22, 22, 'sp12_h_r_20')
// (23, 22, 'sp12_h_r_23')
// (24, 22, 'sp12_h_l_23')

wire n642;
// (12, 23, 'lutff_7/cout')
// (12, 24, 'carry_in')
// (12, 24, 'carry_in_mux')
// (12, 24, 'lutff_0/in_3')

reg io_33_6_0 = 0;
// (12, 23, 'sp12_h_r_0')
// (13, 23, 'sp12_h_r_3')
// (14, 23, 'sp12_h_r_4')
// (15, 23, 'sp12_h_r_7')
// (16, 23, 'sp12_h_r_8')
// (17, 22, 'neigh_op_tnr_2')
// (17, 23, 'neigh_op_rgt_2')
// (17, 23, 'sp12_h_r_11')
// (17, 24, 'neigh_op_bnr_2')
// (18, 22, 'neigh_op_top_2')
// (18, 23, 'lutff_2/out')
// (18, 23, 'sp12_h_r_12')
// (18, 24, 'neigh_op_bot_2')
// (19, 22, 'neigh_op_tnl_2')
// (19, 23, 'neigh_op_lft_2')
// (19, 23, 'sp12_h_r_15')
// (19, 24, 'neigh_op_bnl_2')
// (20, 23, 'sp12_h_r_16')
// (21, 23, 'sp12_h_r_19')
// (22, 23, 'sp12_h_r_20')
// (23, 23, 'sp12_h_r_23')
// (24, 11, 'sp12_h_r_0')
// (24, 11, 'sp12_v_t_23')
// (24, 12, 'sp12_v_b_23')
// (24, 13, 'sp12_v_b_20')
// (24, 14, 'sp12_v_b_19')
// (24, 15, 'sp12_v_b_16')
// (24, 16, 'sp12_v_b_15')
// (24, 17, 'sp12_v_b_12')
// (24, 18, 'sp12_v_b_11')
// (24, 19, 'sp12_v_b_8')
// (24, 20, 'sp12_v_b_7')
// (24, 21, 'sp12_v_b_4')
// (24, 22, 'sp12_v_b_3')
// (24, 23, 'sp12_h_l_23')
// (24, 23, 'sp12_v_b_0')
// (25, 11, 'sp12_h_r_3')
// (25, 11, 'sp4_h_r_3')
// (26, 11, 'sp12_h_r_4')
// (26, 11, 'sp4_h_r_14')
// (27, 11, 'sp12_h_r_7')
// (27, 11, 'sp4_h_r_27')
// (28, 11, 'sp12_h_r_8')
// (28, 11, 'sp4_h_r_38')
// (29, 11, 'sp12_h_r_11')
// (29, 11, 'sp4_h_l_38')
// (29, 11, 'sp4_h_r_6')
// (30, 11, 'sp12_h_r_12')
// (30, 11, 'sp4_h_r_19')
// (31, 11, 'sp12_h_r_15')
// (31, 11, 'sp4_h_r_30')
// (32, 11, 'sp12_h_r_16')
// (32, 11, 'sp4_h_r_43')
// (33, 3, 'span4_vert_t_15')
// (33, 4, 'span4_vert_b_15')
// (33, 5, 'span4_vert_b_11')
// (33, 6, 'io_0/D_OUT_0')
// (33, 6, 'io_0/PAD')
// (33, 6, 'local_g1_7')
// (33, 6, 'span4_vert_b_7')
// (33, 7, 'span4_vert_b_3')
// (33, 7, 'span4_vert_t_15')
// (33, 8, 'span4_vert_b_15')
// (33, 9, 'span4_vert_b_11')
// (33, 10, 'span4_vert_b_7')
// (33, 11, 'span12_horz_16')
// (33, 11, 'span4_horz_43')
// (33, 11, 'span4_vert_b_3')

reg n644 = 0;
// (12, 24, 'sp12_h_r_1')
// (13, 24, 'sp12_h_r_2')
// (14, 24, 'sp12_h_r_5')
// (15, 24, 'sp12_h_r_6')
// (16, 24, 'sp12_h_r_9')
// (17, 24, 'sp12_h_r_10')
// (18, 24, 'local_g0_5')
// (18, 24, 'lutff_1/in_0')
// (18, 24, 'sp12_h_r_13')
// (19, 24, 'sp12_h_r_14')
// (20, 24, 'sp12_h_r_17')
// (21, 24, 'sp12_h_r_18')
// (22, 24, 'sp12_h_r_21')
// (23, 16, 'neigh_op_tnr_7')
// (23, 17, 'neigh_op_rgt_7')
// (23, 18, 'neigh_op_bnr_7')
// (23, 24, 'sp12_h_r_22')
// (24, 12, 'sp12_v_t_22')
// (24, 13, 'sp12_v_b_22')
// (24, 14, 'sp12_v_b_21')
// (24, 15, 'sp12_v_b_18')
// (24, 16, 'neigh_op_top_7')
// (24, 16, 'sp12_v_b_17')
// (24, 17, 'lutff_7/out')
// (24, 17, 'sp12_v_b_14')
// (24, 18, 'neigh_op_bot_7')
// (24, 18, 'sp12_v_b_13')
// (24, 19, 'sp12_v_b_10')
// (24, 20, 'sp12_v_b_9')
// (24, 21, 'sp12_v_b_6')
// (24, 22, 'sp12_v_b_5')
// (24, 23, 'sp12_v_b_2')
// (24, 24, 'sp12_h_l_22')
// (24, 24, 'sp12_v_b_1')
// (25, 16, 'neigh_op_tnl_7')
// (25, 17, 'neigh_op_lft_7')
// (25, 18, 'neigh_op_bnl_7')

wire n645;
// (13, 5, 'sp4_r_v_b_45')
// (13, 6, 'sp4_r_v_b_32')
// (13, 7, 'local_g3_5')
// (13, 7, 'lutff_2/in_0')
// (13, 7, 'sp4_r_v_b_21')
// (13, 8, 'sp4_r_v_b_8')
// (14, 4, 'sp4_v_t_45')
// (14, 5, 'sp4_v_b_45')
// (14, 6, 'sp4_v_b_32')
// (14, 7, 'neigh_op_tnr_7')
// (14, 7, 'sp4_v_b_21')
// (14, 8, 'neigh_op_rgt_7')
// (14, 8, 'sp4_h_r_3')
// (14, 8, 'sp4_v_b_8')
// (14, 9, 'neigh_op_bnr_7')
// (15, 7, 'neigh_op_top_7')
// (15, 8, 'lutff_7/out')
// (15, 8, 'sp4_h_r_14')
// (15, 9, 'neigh_op_bot_7')
// (16, 7, 'neigh_op_tnl_7')
// (16, 8, 'neigh_op_lft_7')
// (16, 8, 'sp4_h_r_27')
// (16, 9, 'neigh_op_bnl_7')
// (17, 8, 'sp4_h_r_38')
// (18, 8, 'sp4_h_l_38')

reg n646 = 0;
// (13, 6, 'neigh_op_tnr_0')
// (13, 7, 'local_g3_0')
// (13, 7, 'lutff_3/in_0')
// (13, 7, 'neigh_op_rgt_0')
// (13, 8, 'neigh_op_bnr_0')
// (14, 6, 'neigh_op_top_0')
// (14, 7, 'local_g1_0')
// (14, 7, 'lutff_0/in_1')
// (14, 7, 'lutff_0/out')
// (14, 8, 'neigh_op_bot_0')
// (15, 6, 'neigh_op_tnl_0')
// (15, 7, 'local_g1_0')
// (15, 7, 'lutff_5/in_2')
// (15, 7, 'neigh_op_lft_0')
// (15, 8, 'neigh_op_bnl_0')

reg n647 = 0;
// (13, 6, 'neigh_op_tnr_1')
// (13, 7, 'local_g2_1')
// (13, 7, 'lutff_2/in_3')
// (13, 7, 'neigh_op_rgt_1')
// (13, 8, 'neigh_op_bnr_1')
// (14, 6, 'neigh_op_top_1')
// (14, 7, 'local_g1_1')
// (14, 7, 'lutff_1/in_1')
// (14, 7, 'lutff_1/out')
// (14, 8, 'neigh_op_bot_1')
// (15, 6, 'neigh_op_tnl_1')
// (15, 7, 'local_g0_1')
// (15, 7, 'local_g1_1')
// (15, 7, 'lutff_1/in_1')
// (15, 7, 'lutff_6/in_1')
// (15, 7, 'neigh_op_lft_1')
// (15, 8, 'local_g2_1')
// (15, 8, 'lutff_1/in_0')
// (15, 8, 'neigh_op_bnl_1')

reg n648 = 0;
// (13, 6, 'neigh_op_tnr_2')
// (13, 7, 'local_g2_2')
// (13, 7, 'lutff_1/in_3')
// (13, 7, 'neigh_op_rgt_2')
// (13, 8, 'local_g0_2')
// (13, 8, 'lutff_6/in_0')
// (13, 8, 'neigh_op_bnr_2')
// (14, 6, 'neigh_op_top_2')
// (14, 7, 'local_g1_2')
// (14, 7, 'lutff_2/in_1')
// (14, 7, 'lutff_2/out')
// (14, 8, 'neigh_op_bot_2')
// (15, 6, 'neigh_op_tnl_2')
// (15, 7, 'local_g1_2')
// (15, 7, 'lutff_1/in_0')
// (15, 7, 'lutff_6/in_3')
// (15, 7, 'neigh_op_lft_2')
// (15, 8, 'local_g2_2')
// (15, 8, 'lutff_0/in_0')
// (15, 8, 'lutff_7/in_3')
// (15, 8, 'neigh_op_bnl_2')

reg n649 = 0;
// (13, 6, 'neigh_op_tnr_3')
// (13, 7, 'neigh_op_rgt_3')
// (13, 8, 'neigh_op_bnr_3')
// (14, 6, 'neigh_op_top_3')
// (14, 7, 'local_g1_3')
// (14, 7, 'lutff_3/in_1')
// (14, 7, 'lutff_3/out')
// (14, 8, 'neigh_op_bot_3')
// (15, 6, 'neigh_op_tnl_3')
// (15, 7, 'local_g1_3')
// (15, 7, 'lutff_5/in_1')
// (15, 7, 'neigh_op_lft_3')
// (15, 8, 'neigh_op_bnl_3')

reg n650 = 0;
// (13, 6, 'neigh_op_tnr_4')
// (13, 7, 'neigh_op_rgt_4')
// (13, 8, 'neigh_op_bnr_4')
// (14, 6, 'neigh_op_top_4')
// (14, 7, 'local_g3_4')
// (14, 7, 'lutff_4/in_1')
// (14, 7, 'lutff_4/out')
// (14, 8, 'neigh_op_bot_4')
// (15, 6, 'neigh_op_tnl_4')
// (15, 7, 'local_g1_4')
// (15, 7, 'lutff_5/in_0')
// (15, 7, 'neigh_op_lft_4')
// (15, 8, 'neigh_op_bnl_4')

reg n651 = 0;
// (13, 6, 'neigh_op_tnr_5')
// (13, 7, 'neigh_op_rgt_5')
// (13, 8, 'neigh_op_bnr_5')
// (14, 6, 'neigh_op_top_5')
// (14, 7, 'local_g3_5')
// (14, 7, 'lutff_5/in_1')
// (14, 7, 'lutff_5/out')
// (14, 8, 'neigh_op_bot_5')
// (15, 6, 'neigh_op_tnl_5')
// (15, 7, 'local_g1_5')
// (15, 7, 'lutff_5/in_3')
// (15, 7, 'neigh_op_lft_5')
// (15, 8, 'neigh_op_bnl_5')

reg n652 = 0;
// (13, 6, 'sp4_r_v_b_40')
// (13, 7, 'local_g1_5')
// (13, 7, 'lutff_1/in_1')
// (13, 7, 'sp4_r_v_b_29')
// (13, 8, 'sp4_r_v_b_16')
// (13, 9, 'sp4_r_v_b_5')
// (14, 5, 'sp4_v_t_40')
// (14, 6, 'sp4_v_b_40')
// (14, 7, 'sp4_v_b_29')
// (14, 8, 'neigh_op_tnr_0')
// (14, 8, 'sp4_v_b_16')
// (14, 9, 'neigh_op_rgt_0')
// (14, 9, 'sp4_h_r_5')
// (14, 9, 'sp4_v_b_5')
// (14, 10, 'neigh_op_bnr_0')
// (15, 8, 'neigh_op_top_0')
// (15, 9, 'lutff_0/out')
// (15, 9, 'sp4_h_r_16')
// (15, 10, 'neigh_op_bot_0')
// (16, 8, 'neigh_op_tnl_0')
// (16, 9, 'neigh_op_lft_0')
// (16, 9, 'sp4_h_r_29')
// (16, 10, 'neigh_op_bnl_0')
// (17, 9, 'sp4_h_r_40')
// (18, 9, 'sp4_h_l_40')

reg n653 = 0;
// (13, 6, 'sp4_r_v_b_42')
// (13, 7, 'sp4_r_v_b_31')
// (13, 8, 'local_g3_2')
// (13, 8, 'lutff_6/in_1')
// (13, 8, 'sp4_r_v_b_18')
// (13, 9, 'sp4_r_v_b_7')
// (14, 5, 'sp4_v_t_42')
// (14, 6, 'sp4_v_b_42')
// (14, 7, 'sp4_v_b_31')
// (14, 8, 'neigh_op_tnr_1')
// (14, 8, 'sp4_v_b_18')
// (14, 9, 'neigh_op_rgt_1')
// (14, 9, 'sp4_h_r_7')
// (14, 9, 'sp4_v_b_7')
// (14, 10, 'neigh_op_bnr_1')
// (15, 8, 'neigh_op_top_1')
// (15, 9, 'lutff_1/out')
// (15, 9, 'sp4_h_r_18')
// (15, 10, 'neigh_op_bot_1')
// (16, 8, 'neigh_op_tnl_1')
// (16, 9, 'neigh_op_lft_1')
// (16, 9, 'sp4_h_r_31')
// (16, 10, 'neigh_op_bnl_1')
// (17, 9, 'sp4_h_r_42')
// (18, 9, 'sp4_h_l_42')

reg n654 = 0;
// (13, 7, 'local_g1_0')
// (13, 7, 'lutff_1/in_0')
// (13, 7, 'sp4_h_r_8')
// (14, 7, 'sp4_h_r_21')
// (15, 7, 'sp4_h_r_32')
// (16, 7, 'sp4_h_r_45')
// (17, 6, 'neigh_op_tnr_0')
// (17, 7, 'neigh_op_rgt_0')
// (17, 7, 'sp4_h_l_45')
// (17, 7, 'sp4_h_r_5')
// (17, 8, 'neigh_op_bnr_0')
// (18, 6, 'neigh_op_top_0')
// (18, 7, 'lutff_0/out')
// (18, 7, 'sp4_h_r_16')
// (18, 8, 'neigh_op_bot_0')
// (19, 6, 'neigh_op_tnl_0')
// (19, 7, 'neigh_op_lft_0')
// (19, 7, 'sp4_h_r_29')
// (19, 8, 'neigh_op_bnl_0')
// (20, 7, 'sp4_h_r_40')
// (21, 7, 'sp4_h_l_40')

wire n655;
// (13, 7, 'lutff_1/lout')
// (13, 7, 'lutff_2/in_2')

wire n656;
// (13, 7, 'lutff_2/lout')
// (13, 7, 'lutff_3/in_2')

wire n657;
// (13, 8, 'neigh_op_tnr_0')
// (13, 9, 'neigh_op_rgt_0')
// (13, 10, 'neigh_op_bnr_0')
// (14, 8, 'neigh_op_top_0')
// (14, 9, 'local_g1_0')
// (14, 9, 'lutff_0/out')
// (14, 9, 'lutff_4/in_3')
// (14, 10, 'neigh_op_bot_0')
// (15, 8, 'neigh_op_tnl_0')
// (15, 9, 'neigh_op_lft_0')
// (15, 10, 'neigh_op_bnl_0')

reg n658 = 0;
// (13, 9, 'neigh_op_tnr_0')
// (13, 10, 'neigh_op_rgt_0')
// (13, 11, 'neigh_op_bnr_0')
// (14, 9, 'neigh_op_top_0')
// (14, 10, 'lutff_0/out')
// (14, 11, 'local_g1_0')
// (14, 11, 'lutff_2/in_3')
// (14, 11, 'neigh_op_bot_0')
// (15, 9, 'neigh_op_tnl_0')
// (15, 10, 'neigh_op_lft_0')
// (15, 11, 'neigh_op_bnl_0')

reg n659 = 0;
// (13, 9, 'neigh_op_tnr_1')
// (13, 10, 'neigh_op_rgt_1')
// (13, 11, 'neigh_op_bnr_1')
// (14, 9, 'neigh_op_top_1')
// (14, 10, 'lutff_1/out')
// (14, 11, 'local_g1_1')
// (14, 11, 'lutff_3/in_3')
// (14, 11, 'neigh_op_bot_1')
// (15, 9, 'neigh_op_tnl_1')
// (15, 10, 'neigh_op_lft_1')
// (15, 11, 'neigh_op_bnl_1')

reg n660 = 0;
// (13, 9, 'neigh_op_tnr_2')
// (13, 10, 'neigh_op_rgt_2')
// (13, 11, 'neigh_op_bnr_2')
// (14, 9, 'neigh_op_top_2')
// (14, 10, 'lutff_2/out')
// (14, 11, 'neigh_op_bot_2')
// (15, 9, 'neigh_op_tnl_2')
// (15, 10, 'neigh_op_lft_2')
// (15, 11, 'local_g2_2')
// (15, 11, 'lutff_1/in_3')
// (15, 11, 'neigh_op_bnl_2')

reg n661 = 0;
// (13, 9, 'neigh_op_tnr_3')
// (13, 10, 'local_g3_3')
// (13, 10, 'lutff_1/in_3')
// (13, 10, 'neigh_op_rgt_3')
// (13, 11, 'neigh_op_bnr_3')
// (14, 9, 'neigh_op_top_3')
// (14, 10, 'lutff_3/out')
// (14, 11, 'neigh_op_bot_3')
// (15, 9, 'neigh_op_tnl_3')
// (15, 10, 'neigh_op_lft_3')
// (15, 11, 'neigh_op_bnl_3')

reg n662 = 0;
// (13, 9, 'neigh_op_tnr_4')
// (13, 10, 'neigh_op_rgt_4')
// (13, 11, 'neigh_op_bnr_4')
// (14, 9, 'neigh_op_top_4')
// (14, 10, 'lutff_4/out')
// (14, 11, 'local_g1_4')
// (14, 11, 'lutff_6/in_3')
// (14, 11, 'neigh_op_bot_4')
// (15, 9, 'neigh_op_tnl_4')
// (15, 10, 'neigh_op_lft_4')
// (15, 11, 'neigh_op_bnl_4')

reg n663 = 0;
// (13, 9, 'neigh_op_tnr_5')
// (13, 10, 'neigh_op_rgt_5')
// (13, 11, 'neigh_op_bnr_5')
// (14, 9, 'neigh_op_top_5')
// (14, 10, 'lutff_5/out')
// (14, 11, 'local_g1_5')
// (14, 11, 'lutff_7/in_3')
// (14, 11, 'neigh_op_bot_5')
// (15, 9, 'neigh_op_tnl_5')
// (15, 10, 'neigh_op_lft_5')
// (15, 11, 'neigh_op_bnl_5')

reg n664 = 0;
// (13, 9, 'neigh_op_tnr_7')
// (13, 10, 'local_g3_7')
// (13, 10, 'lutff_7/in_3')
// (13, 10, 'neigh_op_rgt_7')
// (13, 11, 'neigh_op_bnr_7')
// (14, 9, 'neigh_op_top_7')
// (14, 10, 'lutff_7/out')
// (14, 11, 'neigh_op_bot_7')
// (15, 9, 'neigh_op_tnl_7')
// (15, 10, 'neigh_op_lft_7')
// (15, 11, 'neigh_op_bnl_7')

reg n665 = 0;
// (13, 9, 'sp4_r_v_b_36')
// (13, 10, 'neigh_op_tnr_6')
// (13, 10, 'sp4_r_v_b_25')
// (13, 11, 'neigh_op_rgt_6')
// (13, 11, 'sp4_r_v_b_12')
// (13, 12, 'neigh_op_bnr_6')
// (13, 12, 'sp4_r_v_b_1')
// (14, 8, 'sp4_v_t_36')
// (14, 9, 'local_g2_4')
// (14, 9, 'lutff_3/in_1')
// (14, 9, 'sp4_v_b_36')
// (14, 10, 'neigh_op_top_6')
// (14, 10, 'sp4_v_b_25')
// (14, 11, 'lutff_6/out')
// (14, 11, 'sp4_v_b_12')
// (14, 12, 'neigh_op_bot_6')
// (14, 12, 'sp4_v_b_1')
// (15, 10, 'neigh_op_tnl_6')
// (15, 11, 'neigh_op_lft_6')
// (15, 12, 'neigh_op_bnl_6')

wire n666;
// (13, 9, 'sp4_r_v_b_43')
// (13, 10, 'sp4_r_v_b_30')
// (13, 11, 'neigh_op_tnr_3')
// (13, 11, 'sp4_r_v_b_19')
// (13, 12, 'neigh_op_rgt_3')
// (13, 12, 'sp4_r_v_b_6')
// (13, 13, 'neigh_op_bnr_3')
// (14, 8, 'sp4_v_t_43')
// (14, 9, 'local_g3_3')
// (14, 9, 'lutff_5/in_1')
// (14, 9, 'sp4_v_b_43')
// (14, 10, 'sp4_v_b_30')
// (14, 11, 'neigh_op_top_3')
// (14, 11, 'sp4_v_b_19')
// (14, 12, 'lutff_3/out')
// (14, 12, 'sp4_v_b_6')
// (14, 13, 'neigh_op_bot_3')
// (15, 11, 'neigh_op_tnl_3')
// (15, 12, 'neigh_op_lft_3')
// (15, 13, 'neigh_op_bnl_3')

reg n667 = 0;
// (13, 9, 'sp4_r_v_b_44')
// (13, 10, 'neigh_op_tnr_2')
// (13, 10, 'sp4_r_v_b_33')
// (13, 11, 'neigh_op_rgt_2')
// (13, 11, 'sp4_r_v_b_20')
// (13, 12, 'neigh_op_bnr_2')
// (13, 12, 'sp4_r_v_b_9')
// (14, 8, 'sp4_v_t_44')
// (14, 9, 'local_g3_4')
// (14, 9, 'lutff_0/in_3')
// (14, 9, 'sp4_v_b_44')
// (14, 10, 'neigh_op_top_2')
// (14, 10, 'sp4_v_b_33')
// (14, 11, 'lutff_2/out')
// (14, 11, 'sp4_v_b_20')
// (14, 12, 'neigh_op_bot_2')
// (14, 12, 'sp4_v_b_9')
// (15, 10, 'neigh_op_tnl_2')
// (15, 11, 'neigh_op_lft_2')
// (15, 12, 'neigh_op_bnl_2')

reg n668 = 0;
// (13, 10, 'local_g0_3')
// (13, 10, 'lutff_0/in_3')
// (13, 10, 'sp4_h_r_11')
// (14, 10, 'sp4_h_r_22')
// (15, 9, 'neigh_op_tnr_7')
// (15, 10, 'neigh_op_rgt_7')
// (15, 10, 'sp4_h_r_35')
// (15, 11, 'neigh_op_bnr_7')
// (16, 9, 'neigh_op_top_7')
// (16, 10, 'lutff_7/out')
// (16, 10, 'sp4_h_r_46')
// (16, 11, 'neigh_op_bot_7')
// (17, 9, 'neigh_op_tnl_7')
// (17, 10, 'neigh_op_lft_7')
// (17, 10, 'sp4_h_l_46')
// (17, 11, 'neigh_op_bnl_7')

reg n669 = 0;
// (13, 10, 'local_g0_7')
// (13, 10, 'lutff_4/in_3')
// (13, 10, 'sp4_h_r_7')
// (14, 10, 'sp4_h_r_18')
// (15, 9, 'neigh_op_tnr_5')
// (15, 10, 'neigh_op_rgt_5')
// (15, 10, 'sp4_h_r_31')
// (15, 11, 'neigh_op_bnr_5')
// (16, 9, 'neigh_op_top_5')
// (16, 10, 'lutff_5/out')
// (16, 10, 'sp4_h_r_42')
// (16, 11, 'neigh_op_bot_5')
// (17, 9, 'neigh_op_tnl_5')
// (17, 10, 'neigh_op_lft_5')
// (17, 10, 'sp4_h_l_42')
// (17, 11, 'neigh_op_bnl_5')

reg n670 = 0;
// (13, 10, 'neigh_op_tnr_3')
// (13, 11, 'neigh_op_rgt_3')
// (13, 12, 'neigh_op_bnr_3')
// (14, 10, 'neigh_op_top_3')
// (14, 11, 'lutff_3/out')
// (14, 12, 'local_g1_3')
// (14, 12, 'lutff_0/in_0')
// (14, 12, 'neigh_op_bot_3')
// (15, 10, 'neigh_op_tnl_3')
// (15, 11, 'neigh_op_lft_3')
// (15, 12, 'neigh_op_bnl_3')

reg n671 = 0;
// (13, 10, 'neigh_op_tnr_7')
// (13, 11, 'neigh_op_rgt_7')
// (13, 12, 'neigh_op_bnr_7')
// (14, 10, 'neigh_op_top_7')
// (14, 11, 'lutff_7/out')
// (14, 12, 'local_g0_7')
// (14, 12, 'lutff_0/in_3')
// (14, 12, 'neigh_op_bot_7')
// (15, 10, 'neigh_op_tnl_7')
// (15, 11, 'neigh_op_lft_7')
// (15, 12, 'neigh_op_bnl_7')

reg n672 = 0;
// (13, 10, 'sp4_h_r_2')
// (14, 9, 'neigh_op_tnr_5')
// (14, 9, 'sp4_r_v_b_39')
// (14, 10, 'local_g0_2')
// (14, 10, 'lutff_global/cen')
// (14, 10, 'neigh_op_rgt_5')
// (14, 10, 'sp4_h_r_15')
// (14, 10, 'sp4_r_v_b_26')
// (14, 11, 'neigh_op_bnr_5')
// (14, 11, 'sp4_r_v_b_15')
// (14, 12, 'sp4_r_v_b_2')
// (15, 8, 'sp4_v_t_39')
// (15, 9, 'neigh_op_top_5')
// (15, 9, 'sp4_r_v_b_38')
// (15, 9, 'sp4_v_b_39')
// (15, 10, 'local_g2_5')
// (15, 10, 'lutff_5/in_2')
// (15, 10, 'lutff_5/out')
// (15, 10, 'sp4_h_r_10')
// (15, 10, 'sp4_h_r_26')
// (15, 10, 'sp4_r_v_b_27')
// (15, 10, 'sp4_v_b_26')
// (15, 11, 'neigh_op_bot_5')
// (15, 11, 'sp4_r_v_b_14')
// (15, 11, 'sp4_v_b_15')
// (15, 12, 'sp4_r_v_b_3')
// (15, 12, 'sp4_v_b_2')
// (16, 7, 'sp4_r_v_b_42')
// (16, 8, 'sp4_r_v_b_31')
// (16, 8, 'sp4_v_t_38')
// (16, 9, 'neigh_op_tnl_5')
// (16, 9, 'sp4_r_v_b_18')
// (16, 9, 'sp4_v_b_38')
// (16, 10, 'local_g3_3')
// (16, 10, 'lutff_global/cen')
// (16, 10, 'neigh_op_lft_5')
// (16, 10, 'sp4_h_r_23')
// (16, 10, 'sp4_h_r_39')
// (16, 10, 'sp4_r_v_b_7')
// (16, 10, 'sp4_v_b_27')
// (16, 11, 'neigh_op_bnl_5')
// (16, 11, 'sp4_v_b_14')
// (16, 12, 'sp4_v_b_3')
// (17, 6, 'sp4_v_t_42')
// (17, 7, 'sp4_v_b_42')
// (17, 8, 'sp4_v_b_31')
// (17, 9, 'local_g0_2')
// (17, 9, 'lutff_global/cen')
// (17, 9, 'sp4_v_b_18')
// (17, 10, 'sp4_h_l_39')
// (17, 10, 'sp4_h_r_2')
// (17, 10, 'sp4_h_r_34')
// (17, 10, 'sp4_v_b_7')
// (18, 7, 'sp4_r_v_b_47')
// (18, 8, 'sp4_r_v_b_34')
// (18, 9, 'sp4_r_v_b_23')
// (18, 10, 'sp4_h_r_15')
// (18, 10, 'sp4_h_r_47')
// (18, 10, 'sp4_r_v_b_10')
// (19, 6, 'sp4_v_t_47')
// (19, 7, 'sp4_v_b_47')
// (19, 8, 'local_g2_2')
// (19, 8, 'lutff_global/cen')
// (19, 8, 'sp4_v_b_34')
// (19, 9, 'sp4_v_b_23')
// (19, 10, 'sp4_h_l_47')
// (19, 10, 'sp4_h_r_26')
// (19, 10, 'sp4_v_b_10')
// (20, 10, 'sp4_h_r_39')
// (21, 10, 'sp4_h_l_39')

reg n673 = 0;
// (13, 10, 'sp4_r_v_b_36')
// (13, 11, 'sp4_r_v_b_25')
// (13, 12, 'sp4_r_v_b_12')
// (13, 13, 'sp4_r_v_b_1')
// (13, 14, 'sp4_r_v_b_47')
// (13, 15, 'sp4_r_v_b_34')
// (13, 16, 'neigh_op_tnr_5')
// (13, 16, 'sp4_r_v_b_23')
// (13, 17, 'neigh_op_rgt_5')
// (13, 17, 'sp4_r_v_b_10')
// (13, 18, 'neigh_op_bnr_5')
// (14, 9, 'sp4_v_t_36')
// (14, 10, 'local_g3_4')
// (14, 10, 'lutff_2/in_3')
// (14, 10, 'sp4_v_b_36')
// (14, 11, 'sp4_v_b_25')
// (14, 12, 'sp4_v_b_12')
// (14, 13, 'sp4_v_b_1')
// (14, 13, 'sp4_v_t_47')
// (14, 14, 'sp4_v_b_47')
// (14, 15, 'sp4_v_b_34')
// (14, 16, 'neigh_op_top_5')
// (14, 16, 'sp4_v_b_23')
// (14, 17, 'lutff_5/out')
// (14, 17, 'sp4_v_b_10')
// (14, 18, 'neigh_op_bot_5')
// (15, 16, 'neigh_op_tnl_5')
// (15, 17, 'neigh_op_lft_5')
// (15, 18, 'neigh_op_bnl_5')

wire n674;
// (13, 11, 'lutff_0/lout')
// (13, 11, 'lutff_1/in_2')

wire n675;
// (13, 11, 'lutff_4/lout')
// (13, 11, 'lutff_5/in_2')

wire n676;
// (13, 11, 'neigh_op_tnr_2')
// (13, 12, 'neigh_op_rgt_2')
// (13, 13, 'neigh_op_bnr_2')
// (14, 11, 'neigh_op_top_2')
// (14, 12, 'local_g0_2')
// (14, 12, 'lutff_1/in_3')
// (14, 12, 'lutff_2/out')
// (14, 13, 'neigh_op_bot_2')
// (15, 11, 'neigh_op_tnl_2')
// (15, 12, 'neigh_op_lft_2')
// (15, 13, 'neigh_op_bnl_2')

reg n677 = 0;
// (13, 11, 'sp4_r_v_b_36')
// (13, 12, 'neigh_op_tnr_6')
// (13, 12, 'sp4_r_v_b_25')
// (13, 13, 'neigh_op_rgt_6')
// (13, 13, 'sp4_r_v_b_12')
// (13, 14, 'neigh_op_bnr_6')
// (13, 14, 'sp4_r_v_b_1')
// (14, 10, 'sp4_v_t_36')
// (14, 11, 'sp4_v_b_36')
// (14, 12, 'neigh_op_top_6')
// (14, 12, 'sp4_v_b_25')
// (14, 13, 'lutff_6/out')
// (14, 13, 'sp4_v_b_12')
// (14, 14, 'neigh_op_bot_6')
// (14, 14, 'sp4_h_r_7')
// (14, 14, 'sp4_v_b_1')
// (15, 12, 'neigh_op_tnl_6')
// (15, 13, 'neigh_op_lft_6')
// (15, 14, 'neigh_op_bnl_6')
// (15, 14, 'sp4_h_r_18')
// (16, 14, 'sp4_h_r_31')
// (17, 14, 'sp4_h_r_42')
// (18, 14, 'sp4_h_l_42')
// (18, 14, 'sp4_h_r_10')
// (19, 14, 'local_g0_7')
// (19, 14, 'lutff_6/in_1')
// (19, 14, 'sp4_h_r_23')
// (20, 14, 'sp4_h_r_34')
// (21, 14, 'sp4_h_r_47')
// (22, 14, 'sp4_h_l_47')

wire n678;
// (13, 12, 'lutff_0/cout')
// (13, 12, 'lutff_1/in_3')

wire n679;
// (13, 12, 'lutff_1/cout')
// (13, 12, 'lutff_2/in_3')

wire n680;
// (13, 12, 'lutff_2/cout')
// (13, 12, 'lutff_3/in_3')

wire n681;
// (13, 12, 'lutff_3/cout')
// (13, 12, 'lutff_4/in_3')

wire n682;
// (13, 12, 'lutff_4/cout')
// (13, 12, 'lutff_5/in_3')

reg n683 = 0;
// (13, 12, 'neigh_op_tnr_0')
// (13, 12, 'sp4_r_v_b_45')
// (13, 13, 'neigh_op_rgt_0')
// (13, 13, 'sp4_r_v_b_32')
// (13, 14, 'neigh_op_bnr_0')
// (13, 14, 'sp4_r_v_b_21')
// (13, 15, 'sp4_r_v_b_8')
// (14, 11, 'sp4_v_t_45')
// (14, 12, 'neigh_op_top_0')
// (14, 12, 'sp4_v_b_45')
// (14, 13, 'lutff_0/out')
// (14, 13, 'sp4_v_b_32')
// (14, 14, 'neigh_op_bot_0')
// (14, 14, 'sp4_v_b_21')
// (14, 15, 'sp4_h_r_8')
// (14, 15, 'sp4_v_b_8')
// (15, 12, 'neigh_op_tnl_0')
// (15, 13, 'neigh_op_lft_0')
// (15, 14, 'neigh_op_bnl_0')
// (15, 15, 'sp4_h_r_21')
// (16, 15, 'sp4_h_r_32')
// (17, 15, 'sp4_h_r_45')
// (18, 15, 'local_g1_3')
// (18, 15, 'lutff_5/in_3')
// (18, 15, 'sp4_h_l_45')
// (18, 15, 'sp4_h_r_11')
// (19, 15, 'sp4_h_r_22')
// (20, 15, 'sp4_h_r_35')
// (21, 15, 'sp4_h_r_46')
// (22, 15, 'sp4_h_l_46')

reg n684 = 0;
// (13, 12, 'neigh_op_tnr_2')
// (13, 13, 'neigh_op_rgt_2')
// (13, 14, 'neigh_op_bnr_2')
// (14, 12, 'neigh_op_top_2')
// (14, 13, 'lutff_2/out')
// (14, 13, 'sp4_h_r_4')
// (14, 14, 'neigh_op_bot_2')
// (15, 12, 'neigh_op_tnl_2')
// (15, 13, 'neigh_op_lft_2')
// (15, 13, 'sp4_h_r_17')
// (15, 14, 'neigh_op_bnl_2')
// (16, 13, 'sp4_h_r_28')
// (17, 13, 'sp4_h_r_41')
// (18, 13, 'sp4_h_l_41')
// (18, 13, 'sp4_h_r_0')
// (19, 13, 'sp4_h_r_13')
// (20, 13, 'sp4_h_r_24')
// (21, 13, 'local_g2_5')
// (21, 13, 'lutff_2/in_3')
// (21, 13, 'sp4_h_r_37')
// (22, 13, 'sp4_h_l_37')

reg n685 = 0;
// (13, 12, 'neigh_op_tnr_3')
// (13, 13, 'neigh_op_rgt_3')
// (13, 14, 'neigh_op_bnr_3')
// (14, 4, 'sp12_v_t_22')
// (14, 5, 'sp12_v_b_22')
// (14, 6, 'sp12_v_b_21')
// (14, 7, 'sp12_v_b_18')
// (14, 8, 'sp12_v_b_17')
// (14, 9, 'sp12_v_b_14')
// (14, 10, 'sp12_v_b_13')
// (14, 11, 'sp12_v_b_10')
// (14, 12, 'neigh_op_top_3')
// (14, 12, 'sp12_v_b_9')
// (14, 13, 'lutff_3/out')
// (14, 13, 'sp12_v_b_6')
// (14, 14, 'neigh_op_bot_3')
// (14, 14, 'sp12_v_b_5')
// (14, 15, 'sp12_v_b_2')
// (14, 16, 'sp12_h_r_1')
// (14, 16, 'sp12_v_b_1')
// (15, 12, 'neigh_op_tnl_3')
// (15, 13, 'neigh_op_lft_3')
// (15, 14, 'neigh_op_bnl_3')
// (15, 16, 'sp12_h_r_2')
// (16, 16, 'sp12_h_r_5')
// (17, 16, 'sp12_h_r_6')
// (18, 16, 'sp12_h_r_9')
// (19, 16, 'sp12_h_r_10')
// (20, 16, 'sp12_h_r_13')
// (21, 16, 'local_g1_6')
// (21, 16, 'lutff_6/in_3')
// (21, 16, 'sp12_h_r_14')
// (22, 16, 'sp12_h_r_17')
// (23, 16, 'sp12_h_r_18')
// (24, 16, 'sp12_h_r_21')
// (25, 16, 'sp12_h_r_22')
// (26, 16, 'sp12_h_l_22')

reg n686 = 0;
// (13, 12, 'neigh_op_tnr_4')
// (13, 13, 'neigh_op_rgt_4')
// (13, 14, 'neigh_op_bnr_4')
// (14, 12, 'neigh_op_top_4')
// (14, 13, 'lutff_4/out')
// (14, 13, 'sp4_r_v_b_41')
// (14, 14, 'neigh_op_bot_4')
// (14, 14, 'sp4_r_v_b_28')
// (14, 15, 'sp4_r_v_b_17')
// (14, 16, 'sp4_r_v_b_4')
// (15, 12, 'neigh_op_tnl_4')
// (15, 12, 'sp4_v_t_41')
// (15, 13, 'neigh_op_lft_4')
// (15, 13, 'sp4_v_b_41')
// (15, 14, 'neigh_op_bnl_4')
// (15, 14, 'sp4_v_b_28')
// (15, 15, 'sp4_v_b_17')
// (15, 16, 'sp4_h_r_10')
// (15, 16, 'sp4_v_b_4')
// (16, 16, 'sp4_h_r_23')
// (17, 16, 'sp4_h_r_34')
// (18, 16, 'sp4_h_r_47')
// (19, 16, 'sp4_h_l_47')
// (19, 16, 'sp4_h_r_10')
// (20, 16, 'sp4_h_r_23')
// (21, 16, 'sp4_h_r_34')
// (22, 16, 'local_g2_7')
// (22, 16, 'lutff_4/in_3')
// (22, 16, 'sp4_h_r_47')
// (23, 16, 'sp4_h_l_47')

reg n687 = 0;
// (13, 12, 'neigh_op_tnr_5')
// (13, 13, 'neigh_op_rgt_5')
// (13, 14, 'neigh_op_bnr_5')
// (14, 6, 'sp12_v_t_22')
// (14, 7, 'sp12_v_b_22')
// (14, 8, 'sp12_v_b_21')
// (14, 9, 'sp12_v_b_18')
// (14, 10, 'sp12_v_b_17')
// (14, 11, 'sp12_v_b_14')
// (14, 12, 'neigh_op_top_5')
// (14, 12, 'sp12_v_b_13')
// (14, 13, 'lutff_5/out')
// (14, 13, 'sp12_v_b_10')
// (14, 14, 'neigh_op_bot_5')
// (14, 14, 'sp12_v_b_9')
// (14, 15, 'sp12_v_b_6')
// (14, 16, 'sp12_v_b_5')
// (14, 17, 'sp12_v_b_2')
// (14, 18, 'sp12_h_r_1')
// (14, 18, 'sp12_v_b_1')
// (15, 12, 'neigh_op_tnl_5')
// (15, 13, 'neigh_op_lft_5')
// (15, 14, 'neigh_op_bnl_5')
// (15, 18, 'sp12_h_r_2')
// (16, 18, 'sp12_h_r_5')
// (17, 18, 'sp12_h_r_6')
// (18, 18, 'sp12_h_r_9')
// (19, 18, 'local_g1_2')
// (19, 18, 'lutff_6/in_1')
// (19, 18, 'sp12_h_r_10')
// (20, 18, 'sp12_h_r_13')
// (21, 18, 'sp12_h_r_14')
// (22, 18, 'sp12_h_r_17')
// (23, 18, 'sp12_h_r_18')
// (24, 18, 'sp12_h_r_21')
// (25, 18, 'sp12_h_r_22')
// (26, 18, 'sp12_h_l_22')

wire n688;
// (13, 12, 'sp4_r_v_b_46')
// (13, 13, 'sp4_r_v_b_35')
// (13, 14, 'sp4_r_v_b_22')
// (13, 15, 'sp4_r_v_b_11')
// (14, 11, 'sp4_v_t_46')
// (14, 12, 'sp4_v_b_46')
// (14, 13, 'sp4_v_b_35')
// (14, 14, 'sp4_v_b_22')
// (14, 15, 'local_g1_3')
// (14, 15, 'lutff_global/cen')
// (14, 15, 'sp4_h_r_6')
// (14, 15, 'sp4_v_b_11')
// (15, 14, 'neigh_op_tnr_7')
// (15, 15, 'neigh_op_rgt_7')
// (15, 15, 'sp4_h_r_19')
// (15, 16, 'neigh_op_bnr_7')
// (16, 14, 'neigh_op_top_7')
// (16, 15, 'lutff_7/out')
// (16, 15, 'sp4_h_r_30')
// (16, 16, 'neigh_op_bot_7')
// (17, 14, 'neigh_op_tnl_7')
// (17, 15, 'neigh_op_lft_7')
// (17, 15, 'sp4_h_r_43')
// (17, 16, 'neigh_op_bnl_7')
// (17, 16, 'sp4_r_v_b_46')
// (17, 17, 'sp4_r_v_b_35')
// (17, 18, 'sp4_r_v_b_22')
// (17, 19, 'sp4_r_v_b_11')
// (17, 20, 'sp4_r_v_b_39')
// (17, 20, 'sp4_r_v_b_42')
// (17, 21, 'sp4_r_v_b_26')
// (17, 21, 'sp4_r_v_b_31')
// (17, 22, 'sp4_r_v_b_15')
// (17, 22, 'sp4_r_v_b_18')
// (17, 23, 'sp4_r_v_b_2')
// (17, 23, 'sp4_r_v_b_7')
// (18, 15, 'sp4_h_l_43')
// (18, 15, 'sp4_v_t_46')
// (18, 16, 'sp4_v_b_46')
// (18, 17, 'sp4_v_b_35')
// (18, 18, 'sp4_v_b_22')
// (18, 19, 'sp4_v_b_11')
// (18, 19, 'sp4_v_t_39')
// (18, 19, 'sp4_v_t_42')
// (18, 20, 'sp4_v_b_39')
// (18, 20, 'sp4_v_b_42')
// (18, 21, 'sp4_v_b_26')
// (18, 21, 'sp4_v_b_31')
// (18, 22, 'sp4_v_b_15')
// (18, 22, 'sp4_v_b_18')
// (18, 23, 'sp4_h_r_1')
// (18, 23, 'sp4_h_r_2')
// (18, 23, 'sp4_v_b_2')
// (18, 23, 'sp4_v_b_7')
// (19, 23, 'sp4_h_r_12')
// (19, 23, 'sp4_h_r_15')
// (20, 23, 'local_g2_2')
// (20, 23, 'lutff_global/cen')
// (20, 23, 'sp4_h_r_25')
// (20, 23, 'sp4_h_r_26')
// (21, 23, 'sp4_h_r_36')
// (21, 23, 'sp4_h_r_39')
// (21, 24, 'local_g3_3')
// (21, 24, 'lutff_global/cen')
// (21, 24, 'sp4_r_v_b_43')
// (21, 25, 'sp4_r_v_b_30')
// (21, 26, 'sp4_r_v_b_19')
// (21, 27, 'sp4_r_v_b_6')
// (22, 23, 'sp4_h_l_36')
// (22, 23, 'sp4_h_l_39')
// (22, 23, 'sp4_v_t_43')
// (22, 24, 'sp4_v_b_43')
// (22, 25, 'sp4_v_b_30')
// (22, 26, 'sp4_v_b_19')
// (22, 27, 'sp4_v_b_6')

reg n689 = 0;
// (13, 13, 'neigh_op_tnr_0')
// (13, 13, 'sp4_r_v_b_45')
// (13, 14, 'neigh_op_rgt_0')
// (13, 14, 'sp4_r_v_b_32')
// (13, 15, 'neigh_op_bnr_0')
// (13, 15, 'sp4_r_v_b_21')
// (13, 16, 'sp4_r_v_b_8')
// (14, 12, 'sp4_h_r_8')
// (14, 12, 'sp4_v_t_45')
// (14, 13, 'neigh_op_top_0')
// (14, 13, 'sp4_v_b_45')
// (14, 14, 'lutff_0/out')
// (14, 14, 'sp4_v_b_32')
// (14, 15, 'neigh_op_bot_0')
// (14, 15, 'sp4_v_b_21')
// (14, 16, 'sp4_v_b_8')
// (15, 12, 'sp4_h_r_21')
// (15, 13, 'local_g2_0')
// (15, 13, 'lutff_1/in_1')
// (15, 13, 'lutff_4/in_2')
// (15, 13, 'neigh_op_tnl_0')
// (15, 14, 'local_g1_0')
// (15, 14, 'lutff_7/in_0')
// (15, 14, 'neigh_op_lft_0')
// (15, 15, 'neigh_op_bnl_0')
// (16, 12, 'local_g2_0')
// (16, 12, 'lutff_2/in_2')
// (16, 12, 'sp4_h_r_32')
// (17, 12, 'sp4_h_r_45')
// (18, 12, 'sp4_h_l_45')

wire n690;
// (13, 13, 'sp4_h_r_6')
// (14, 13, 'local_g1_3')
// (14, 13, 'lutff_global/cen')
// (14, 13, 'sp4_h_r_19')
// (15, 12, 'neigh_op_tnr_0')
// (15, 13, 'neigh_op_rgt_0')
// (15, 13, 'sp4_h_r_30')
// (15, 14, 'neigh_op_bnr_0')
// (16, 10, 'sp4_r_v_b_36')
// (16, 11, 'sp4_r_v_b_25')
// (16, 12, 'neigh_op_top_0')
// (16, 12, 'sp4_r_v_b_12')
// (16, 13, 'lutff_0/out')
// (16, 13, 'sp4_h_r_43')
// (16, 13, 'sp4_r_v_b_1')
// (16, 14, 'neigh_op_bot_0')
// (17, 9, 'sp4_v_t_36')
// (17, 10, 'sp4_v_b_36')
// (17, 11, 'sp4_v_b_25')
// (17, 12, 'neigh_op_tnl_0')
// (17, 12, 'sp4_v_b_12')
// (17, 13, 'neigh_op_lft_0')
// (17, 13, 'sp4_h_l_43')
// (17, 13, 'sp4_v_b_1')
// (17, 14, 'neigh_op_bnl_0')

wire n691;
// (13, 13, 'sp4_r_v_b_38')
// (13, 14, 'neigh_op_tnr_7')
// (13, 14, 'sp4_r_v_b_27')
// (13, 15, 'neigh_op_rgt_7')
// (13, 15, 'sp4_r_v_b_14')
// (13, 16, 'neigh_op_bnr_7')
// (13, 16, 'sp4_r_v_b_3')
// (14, 12, 'sp4_h_r_3')
// (14, 12, 'sp4_v_t_38')
// (14, 13, 'sp4_v_b_38')
// (14, 14, 'neigh_op_top_7')
// (14, 14, 'sp4_v_b_27')
// (14, 15, 'lutff_7/out')
// (14, 15, 'sp4_v_b_14')
// (14, 16, 'neigh_op_bot_7')
// (14, 16, 'sp4_v_b_3')
// (15, 12, 'local_g1_6')
// (15, 12, 'lutff_1/in_2')
// (15, 12, 'sp4_h_r_14')
// (15, 14, 'neigh_op_tnl_7')
// (15, 15, 'neigh_op_lft_7')
// (15, 16, 'neigh_op_bnl_7')
// (16, 12, 'sp4_h_r_27')
// (17, 12, 'sp4_h_r_38')
// (18, 12, 'sp4_h_l_38')

wire n692;
// (13, 14, 'neigh_op_tnr_0')
// (13, 15, 'neigh_op_rgt_0')
// (13, 16, 'neigh_op_bnr_0')
// (14, 11, 'sp12_v_t_23')
// (14, 12, 'sp12_v_b_23')
// (14, 13, 'sp12_v_b_20')
// (14, 14, 'neigh_op_top_0')
// (14, 14, 'sp12_v_b_19')
// (14, 15, 'lutff_0/out')
// (14, 15, 'sp12_v_b_16')
// (14, 16, 'neigh_op_bot_0')
// (14, 16, 'sp12_v_b_15')
// (14, 17, 'sp12_v_b_12')
// (14, 18, 'sp12_v_b_11')
// (14, 19, 'sp12_v_b_8')
// (14, 20, 'sp12_v_b_7')
// (14, 21, 'sp12_v_b_4')
// (14, 22, 'sp12_v_b_3')
// (14, 23, 'sp12_h_r_0')
// (14, 23, 'sp12_v_b_0')
// (15, 14, 'neigh_op_tnl_0')
// (15, 15, 'neigh_op_lft_0')
// (15, 16, 'neigh_op_bnl_0')
// (15, 23, 'sp12_h_r_3')
// (16, 23, 'sp12_h_r_4')
// (17, 23, 'sp12_h_r_7')
// (18, 23, 'sp12_h_r_8')
// (19, 23, 'sp12_h_r_11')
// (20, 23, 'local_g0_4')
// (20, 23, 'lutff_0/in_2')
// (20, 23, 'sp12_h_r_12')
// (21, 23, 'sp12_h_r_15')
// (22, 23, 'sp12_h_r_16')
// (23, 23, 'sp12_h_r_19')
// (24, 23, 'sp12_h_r_20')
// (25, 23, 'sp12_h_r_23')
// (26, 23, 'sp12_h_l_23')

reg n693 = 0;
// (13, 14, 'neigh_op_tnr_1')
// (13, 15, 'neigh_op_rgt_1')
// (13, 16, 'neigh_op_bnr_1')
// (14, 14, 'neigh_op_top_1')
// (14, 15, 'local_g3_1')
// (14, 15, 'lutff_0/in_0')
// (14, 15, 'lutff_1/out')
// (14, 16, 'neigh_op_bot_1')
// (15, 14, 'neigh_op_tnl_1')
// (15, 15, 'neigh_op_lft_1')
// (15, 16, 'neigh_op_bnl_1')

reg n694 = 0;
// (13, 14, 'neigh_op_tnr_4')
// (13, 15, 'neigh_op_rgt_4')
// (13, 16, 'neigh_op_bnr_4')
// (14, 14, 'neigh_op_top_4')
// (14, 15, 'local_g0_4')
// (14, 15, 'lutff_0/in_2')
// (14, 15, 'lutff_4/out')
// (14, 16, 'neigh_op_bot_4')
// (15, 14, 'neigh_op_tnl_4')
// (15, 15, 'neigh_op_lft_4')
// (15, 16, 'neigh_op_bnl_4')

reg n695 = 0;
// (13, 14, 'sp12_h_r_1')
// (14, 14, 'sp12_h_r_2')
// (15, 14, 'sp12_h_r_5')
// (16, 14, 'sp12_h_r_6')
// (17, 14, 'local_g0_1')
// (17, 14, 'lutff_6/in_1')
// (17, 14, 'sp12_h_r_9')
// (18, 14, 'sp12_h_r_10')
// (19, 14, 'sp12_h_r_13')
// (20, 14, 'sp12_h_r_14')
// (21, 14, 'sp12_h_r_17')
// (22, 14, 'sp12_h_r_18')
// (23, 13, 'neigh_op_tnr_7')
// (23, 14, 'neigh_op_rgt_7')
// (23, 14, 'sp12_h_r_21')
// (23, 15, 'neigh_op_bnr_7')
// (24, 13, 'neigh_op_top_7')
// (24, 14, 'lutff_7/out')
// (24, 14, 'sp12_h_r_22')
// (24, 15, 'neigh_op_bot_7')
// (25, 13, 'neigh_op_tnl_7')
// (25, 14, 'neigh_op_lft_7')
// (25, 14, 'sp12_h_l_22')
// (25, 15, 'neigh_op_bnl_7')

reg n696 = 0;
// (13, 15, 'local_g3_6')
// (13, 15, 'lutff_2/in_3')
// (13, 15, 'neigh_op_tnr_6')
// (13, 16, 'neigh_op_rgt_6')
// (13, 17, 'neigh_op_bnr_6')
// (14, 15, 'local_g0_6')
// (14, 15, 'lutff_5/in_3')
// (14, 15, 'neigh_op_top_6')
// (14, 16, 'local_g3_6')
// (14, 16, 'lutff_0/in_3')
// (14, 16, 'lutff_3/in_0')
// (14, 16, 'lutff_6/in_3')
// (14, 16, 'lutff_6/out')
// (14, 17, 'neigh_op_bot_6')
// (15, 15, 'neigh_op_tnl_6')
// (15, 16, 'neigh_op_lft_6')
// (15, 17, 'neigh_op_bnl_6')

wire n697;
// (13, 15, 'neigh_op_tnr_0')
// (13, 15, 'sp4_r_v_b_45')
// (13, 16, 'neigh_op_rgt_0')
// (13, 16, 'sp4_r_v_b_32')
// (13, 17, 'neigh_op_bnr_0')
// (13, 17, 'sp4_r_v_b_21')
// (13, 18, 'sp4_r_v_b_8')
// (13, 19, 'sp4_r_v_b_46')
// (13, 20, 'sp4_r_v_b_35')
// (13, 21, 'sp4_r_v_b_22')
// (13, 22, 'sp4_r_v_b_11')
// (14, 14, 'sp4_v_t_45')
// (14, 15, 'neigh_op_top_0')
// (14, 15, 'sp4_v_b_45')
// (14, 16, 'lutff_0/out')
// (14, 16, 'sp4_v_b_32')
// (14, 17, 'neigh_op_bot_0')
// (14, 17, 'sp4_v_b_21')
// (14, 18, 'sp4_v_b_8')
// (14, 18, 'sp4_v_t_46')
// (14, 19, 'sp4_v_b_46')
// (14, 20, 'sp4_v_b_35')
// (14, 21, 'sp4_v_b_22')
// (14, 22, 'sp4_h_r_5')
// (14, 22, 'sp4_v_b_11')
// (15, 15, 'neigh_op_tnl_0')
// (15, 16, 'neigh_op_lft_0')
// (15, 17, 'neigh_op_bnl_0')
// (15, 22, 'sp4_h_r_16')
// (16, 22, 'sp4_h_r_29')
// (17, 22, 'sp4_h_r_40')
// (17, 23, 'sp4_r_v_b_40')
// (17, 24, 'sp4_r_v_b_29')
// (17, 25, 'sp4_r_v_b_16')
// (17, 26, 'sp4_r_v_b_5')
// (18, 22, 'local_g0_0')
// (18, 22, 'lutff_0/in_2')
// (18, 22, 'lutff_3/in_1')
// (18, 22, 'lutff_4/in_0')
// (18, 22, 'sp4_h_l_40')
// (18, 22, 'sp4_h_r_5')
// (18, 22, 'sp4_h_r_8')
// (18, 22, 'sp4_v_t_40')
// (18, 23, 'sp4_v_b_40')
// (18, 24, 'sp4_v_b_29')
// (18, 25, 'sp4_v_b_16')
// (18, 26, 'local_g0_5')
// (18, 26, 'lutff_0/in_1')
// (18, 26, 'sp4_v_b_5')
// (19, 22, 'sp4_h_r_16')
// (19, 22, 'sp4_h_r_21')
// (20, 22, 'local_g3_5')
// (20, 22, 'lutff_1/in_3')
// (20, 22, 'lutff_5/in_1')
// (20, 22, 'sp4_h_r_29')
// (20, 22, 'sp4_h_r_32')
// (21, 22, 'sp4_h_r_40')
// (21, 22, 'sp4_h_r_45')
// (22, 22, 'sp4_h_l_40')
// (22, 22, 'sp4_h_l_45')

reg n698 = 0;
// (13, 15, 'neigh_op_tnr_1')
// (13, 16, 'neigh_op_rgt_1')
// (13, 17, 'neigh_op_bnr_1')
// (14, 15, 'neigh_op_top_1')
// (14, 16, 'local_g3_1')
// (14, 16, 'lutff_0/in_2')
// (14, 16, 'lutff_1/out')
// (14, 17, 'neigh_op_bot_1')
// (15, 15, 'neigh_op_tnl_1')
// (15, 16, 'neigh_op_lft_1')
// (15, 17, 'neigh_op_bnl_1')

reg n699 = 0;
// (13, 15, 'neigh_op_tnr_2')
// (13, 16, 'neigh_op_rgt_2')
// (13, 17, 'neigh_op_bnr_2')
// (14, 15, 'neigh_op_top_2')
// (14, 16, 'local_g0_2')
// (14, 16, 'lutff_0/in_0')
// (14, 16, 'lutff_1/in_3')
// (14, 16, 'lutff_2/out')
// (14, 17, 'neigh_op_bot_2')
// (15, 15, 'neigh_op_tnl_2')
// (15, 16, 'neigh_op_lft_2')
// (15, 17, 'neigh_op_bnl_2')

reg n700 = 0;
// (13, 15, 'neigh_op_tnr_3')
// (13, 16, 'neigh_op_rgt_3')
// (13, 17, 'neigh_op_bnr_3')
// (14, 15, 'neigh_op_top_3')
// (14, 16, 'local_g2_3')
// (14, 16, 'lutff_0/in_1')
// (14, 16, 'lutff_2/in_3')
// (14, 16, 'lutff_3/out')
// (14, 17, 'neigh_op_bot_3')
// (15, 15, 'neigh_op_tnl_3')
// (15, 16, 'neigh_op_lft_3')
// (15, 17, 'neigh_op_bnl_3')

reg n701 = 0;
// (13, 15, 'neigh_op_tnr_7')
// (13, 16, 'neigh_op_rgt_7')
// (13, 17, 'neigh_op_bnr_7')
// (14, 15, 'neigh_op_top_7')
// (14, 16, 'local_g2_7')
// (14, 16, 'lutff_4/in_1')
// (14, 16, 'lutff_7/out')
// (14, 17, 'neigh_op_bot_7')
// (15, 15, 'neigh_op_tnl_7')
// (15, 16, 'neigh_op_lft_7')
// (15, 17, 'neigh_op_bnl_7')

wire n702;
// (13, 15, 'sp4_h_r_1')
// (14, 15, 'sp4_h_r_12')
// (15, 14, 'neigh_op_tnr_2')
// (15, 15, 'neigh_op_rgt_2')
// (15, 15, 'sp4_h_r_25')
// (15, 16, 'neigh_op_bnr_2')
// (16, 14, 'neigh_op_top_2')
// (16, 15, 'lutff_2/out')
// (16, 15, 'sp4_h_r_36')
// (16, 16, 'neigh_op_bot_2')
// (16, 16, 'sp4_r_v_b_47')
// (16, 17, 'local_g2_2')
// (16, 17, 'lutff_global/cen')
// (16, 17, 'sp4_r_v_b_34')
// (16, 18, 'sp4_r_v_b_23')
// (16, 19, 'sp4_r_v_b_10')
// (17, 14, 'neigh_op_tnl_2')
// (17, 15, 'neigh_op_lft_2')
// (17, 15, 'sp4_h_l_36')
// (17, 15, 'sp4_h_r_4')
// (17, 15, 'sp4_v_t_47')
// (17, 16, 'neigh_op_bnl_2')
// (17, 16, 'sp4_v_b_47')
// (17, 17, 'sp4_v_b_34')
// (17, 18, 'sp4_v_b_23')
// (17, 19, 'sp4_v_b_10')
// (18, 15, 'sp4_h_r_17')
// (19, 15, 'sp4_h_r_28')
// (20, 15, 'sp4_h_r_41')
// (21, 15, 'sp4_h_l_41')

wire n703;
// (13, 15, 'sp4_h_r_10')
// (14, 15, 'local_g0_7')
// (14, 15, 'lutff_7/in_2')
// (14, 15, 'sp4_h_r_23')
// (15, 11, 'neigh_op_tnr_7')
// (15, 12, 'neigh_op_rgt_7')
// (15, 13, 'neigh_op_bnr_7')
// (15, 15, 'sp4_h_r_34')
// (16, 11, 'neigh_op_top_7')
// (16, 12, 'lutff_7/out')
// (16, 12, 'sp4_r_v_b_47')
// (16, 13, 'neigh_op_bot_7')
// (16, 13, 'sp4_r_v_b_34')
// (16, 14, 'sp4_r_v_b_23')
// (16, 15, 'sp4_h_r_47')
// (16, 15, 'sp4_r_v_b_10')
// (17, 11, 'neigh_op_tnl_7')
// (17, 11, 'sp4_v_t_47')
// (17, 12, 'neigh_op_lft_7')
// (17, 12, 'sp4_v_b_47')
// (17, 13, 'neigh_op_bnl_7')
// (17, 13, 'sp4_v_b_34')
// (17, 14, 'sp4_v_b_23')
// (17, 15, 'sp4_h_l_47')
// (17, 15, 'sp4_h_r_10')
// (17, 15, 'sp4_v_b_10')
// (18, 15, 'sp4_h_r_23')
// (19, 15, 'sp4_h_r_34')
// (20, 15, 'sp4_h_r_47')
// (20, 16, 'sp4_r_v_b_47')
// (20, 17, 'sp4_r_v_b_34')
// (20, 18, 'local_g3_7')
// (20, 18, 'lutff_2/in_0')
// (20, 18, 'sp4_r_v_b_23')
// (20, 19, 'sp4_r_v_b_10')
// (21, 15, 'sp4_h_l_47')
// (21, 15, 'sp4_v_t_47')
// (21, 16, 'sp4_v_b_47')
// (21, 17, 'sp4_v_b_34')
// (21, 18, 'sp4_v_b_23')
// (21, 19, 'sp4_v_b_10')

wire n704;
// (13, 15, 'sp4_r_v_b_39')
// (13, 16, 'sp4_r_v_b_26')
// (13, 17, 'sp4_r_v_b_15')
// (13, 18, 'sp4_r_v_b_2')
// (13, 19, 'sp4_r_v_b_47')
// (13, 20, 'sp4_r_v_b_34')
// (13, 21, 'sp4_r_v_b_23')
// (13, 22, 'sp4_r_v_b_10')
// (14, 14, 'sp4_h_r_8')
// (14, 14, 'sp4_v_t_39')
// (14, 15, 'sp4_v_b_39')
// (14, 16, 'sp4_v_b_26')
// (14, 17, 'sp4_v_b_15')
// (14, 18, 'sp4_v_b_2')
// (14, 18, 'sp4_v_t_47')
// (14, 19, 'sp4_v_b_47')
// (14, 20, 'sp4_v_b_34')
// (14, 21, 'sp4_v_b_23')
// (14, 22, 'local_g0_2')
// (14, 22, 'lutff_global/cen')
// (14, 22, 'sp4_v_b_10')
// (15, 13, 'neigh_op_tnr_0')
// (15, 14, 'neigh_op_rgt_0')
// (15, 14, 'sp4_h_r_21')
// (15, 15, 'neigh_op_bnr_0')
// (16, 13, 'neigh_op_top_0')
// (16, 13, 'sp4_r_v_b_44')
// (16, 14, 'lutff_0/out')
// (16, 14, 'sp4_h_r_32')
// (16, 14, 'sp4_r_v_b_33')
// (16, 15, 'neigh_op_bot_0')
// (16, 15, 'sp4_r_v_b_20')
// (16, 16, 'sp4_r_v_b_9')
// (16, 17, 'sp4_r_v_b_37')
// (16, 18, 'sp4_r_v_b_24')
// (16, 19, 'sp4_r_v_b_13')
// (16, 20, 'sp4_r_v_b_0')
// (16, 21, 'sp4_r_v_b_38')
// (16, 22, 'sp4_r_v_b_27')
// (16, 23, 'sp4_r_v_b_14')
// (16, 24, 'sp4_r_v_b_3')
// (16, 25, 'sp4_r_v_b_38')
// (16, 26, 'local_g1_3')
// (16, 26, 'lutff_global/cen')
// (16, 26, 'sp4_r_v_b_27')
// (16, 27, 'sp4_r_v_b_14')
// (16, 28, 'sp4_r_v_b_3')
// (17, 12, 'sp4_v_t_44')
// (17, 13, 'neigh_op_tnl_0')
// (17, 13, 'sp4_v_b_44')
// (17, 14, 'neigh_op_lft_0')
// (17, 14, 'sp4_h_r_45')
// (17, 14, 'sp4_v_b_33')
// (17, 15, 'neigh_op_bnl_0')
// (17, 15, 'sp4_v_b_20')
// (17, 16, 'sp4_v_b_9')
// (17, 16, 'sp4_v_t_37')
// (17, 17, 'sp4_v_b_37')
// (17, 18, 'sp4_v_b_24')
// (17, 19, 'sp4_v_b_13')
// (17, 20, 'sp4_h_r_6')
// (17, 20, 'sp4_v_b_0')
// (17, 20, 'sp4_v_t_38')
// (17, 21, 'sp4_v_b_38')
// (17, 22, 'sp4_v_b_27')
// (17, 23, 'sp4_v_b_14')
// (17, 24, 'sp4_v_b_3')
// (17, 24, 'sp4_v_t_38')
// (17, 25, 'sp4_v_b_38')
// (17, 26, 'sp4_v_b_27')
// (17, 27, 'sp4_v_b_14')
// (17, 28, 'sp4_v_b_3')
// (18, 14, 'sp4_h_l_45')
// (18, 20, 'local_g1_3')
// (18, 20, 'lutff_global/cen')
// (18, 20, 'sp4_h_r_19')
// (19, 20, 'sp4_h_r_30')
// (20, 20, 'sp4_h_r_43')
// (20, 21, 'sp4_r_v_b_43')
// (20, 22, 'sp4_r_v_b_30')
// (20, 23, 'sp4_r_v_b_19')
// (20, 24, 'sp4_r_v_b_6')
// (21, 20, 'sp4_h_l_43')
// (21, 20, 'sp4_v_t_43')
// (21, 21, 'local_g3_3')
// (21, 21, 'lutff_global/cen')
// (21, 21, 'sp4_v_b_43')
// (21, 22, 'sp4_v_b_30')
// (21, 23, 'sp4_v_b_19')
// (21, 24, 'sp4_v_b_6')

reg n705 = 0;
// (13, 15, 'sp4_r_v_b_43')
// (13, 16, 'sp4_r_v_b_30')
// (13, 17, 'sp4_r_v_b_19')
// (13, 18, 'sp4_r_v_b_6')
// (14, 14, 'sp4_h_r_11')
// (14, 14, 'sp4_v_t_43')
// (14, 15, 'sp4_v_b_43')
// (14, 16, 'sp4_v_b_30')
// (14, 17, 'local_g0_3')
// (14, 17, 'local_g1_3')
// (14, 17, 'lutff_3/in_2')
// (14, 17, 'lutff_4/in_0')
// (14, 17, 'sp4_v_b_19')
// (14, 18, 'sp4_h_r_6')
// (14, 18, 'sp4_v_b_6')
// (15, 14, 'sp4_h_r_22')
// (15, 18, 'sp4_h_r_19')
// (16, 14, 'sp4_h_r_35')
// (16, 18, 'sp4_h_r_30')
// (17, 14, 'sp4_h_r_46')
// (17, 14, 'sp4_r_v_b_46')
// (17, 15, 'neigh_op_tnr_3')
// (17, 15, 'sp4_r_v_b_35')
// (17, 15, 'sp4_r_v_b_38')
// (17, 16, 'neigh_op_rgt_3')
// (17, 16, 'sp4_r_v_b_22')
// (17, 16, 'sp4_r_v_b_27')
// (17, 16, 'sp4_r_v_b_38')
// (17, 17, 'local_g2_3')
// (17, 17, 'lutff_6/in_1')
// (17, 17, 'neigh_op_bnr_3')
// (17, 17, 'sp4_r_v_b_11')
// (17, 17, 'sp4_r_v_b_14')
// (17, 17, 'sp4_r_v_b_27')
// (17, 18, 'sp4_h_r_43')
// (17, 18, 'sp4_r_v_b_14')
// (17, 18, 'sp4_r_v_b_3')
// (17, 19, 'sp4_r_v_b_3')
// (18, 7, 'sp12_v_t_22')
// (18, 8, 'sp12_v_b_22')
// (18, 9, 'sp12_v_b_21')
// (18, 10, 'sp12_v_b_18')
// (18, 11, 'sp12_v_b_17')
// (18, 12, 'sp12_v_b_14')
// (18, 13, 'local_g0_4')
// (18, 13, 'lutff_0/in_2')
// (18, 13, 'lutff_4/in_0')
// (18, 13, 'sp12_v_b_13')
// (18, 13, 'sp4_h_r_4')
// (18, 13, 'sp4_r_v_b_42')
// (18, 13, 'sp4_v_t_46')
// (18, 14, 'local_g0_7')
// (18, 14, 'local_g3_7')
// (18, 14, 'lutff_0/in_2')
// (18, 14, 'lutff_1/in_0')
// (18, 14, 'sp12_v_b_10')
// (18, 14, 'sp4_h_l_46')
// (18, 14, 'sp4_h_r_2')
// (18, 14, 'sp4_h_r_8')
// (18, 14, 'sp4_r_v_b_31')
// (18, 14, 'sp4_r_v_b_47')
// (18, 14, 'sp4_v_b_46')
// (18, 14, 'sp4_v_t_38')
// (18, 15, 'neigh_op_top_3')
// (18, 15, 'sp12_v_b_9')
// (18, 15, 'sp4_r_v_b_18')
// (18, 15, 'sp4_r_v_b_34')
// (18, 15, 'sp4_v_b_35')
// (18, 15, 'sp4_v_b_38')
// (18, 15, 'sp4_v_t_38')
// (18, 16, 'local_g1_3')
// (18, 16, 'lutff_3/in_1')
// (18, 16, 'lutff_3/out')
// (18, 16, 'sp12_v_b_6')
// (18, 16, 'sp4_r_v_b_23')
// (18, 16, 'sp4_r_v_b_7')
// (18, 16, 'sp4_v_b_22')
// (18, 16, 'sp4_v_b_27')
// (18, 16, 'sp4_v_b_38')
// (18, 17, 'neigh_op_bot_3')
// (18, 17, 'sp12_v_b_5')
// (18, 17, 'sp4_r_v_b_10')
// (18, 17, 'sp4_v_b_11')
// (18, 17, 'sp4_v_b_14')
// (18, 17, 'sp4_v_b_27')
// (18, 18, 'sp12_v_b_2')
// (18, 18, 'sp4_h_l_43')
// (18, 18, 'sp4_h_r_3')
// (18, 18, 'sp4_v_b_14')
// (18, 18, 'sp4_v_b_3')
// (18, 19, 'sp12_v_b_1')
// (18, 19, 'sp4_h_r_3')
// (18, 19, 'sp4_v_b_3')
// (19, 12, 'sp4_v_t_42')
// (19, 13, 'sp4_h_r_17')
// (19, 13, 'sp4_v_b_42')
// (19, 13, 'sp4_v_t_47')
// (19, 14, 'sp4_h_r_15')
// (19, 14, 'sp4_h_r_21')
// (19, 14, 'sp4_v_b_31')
// (19, 14, 'sp4_v_b_47')
// (19, 15, 'neigh_op_tnl_3')
// (19, 15, 'sp4_v_b_18')
// (19, 15, 'sp4_v_b_34')
// (19, 16, 'neigh_op_lft_3')
// (19, 16, 'sp4_v_b_23')
// (19, 16, 'sp4_v_b_7')
// (19, 17, 'local_g2_3')
// (19, 17, 'lutff_1/in_0')
// (19, 17, 'lutff_6/in_1')
// (19, 17, 'neigh_op_bnl_3')
// (19, 17, 'sp4_v_b_10')
// (19, 18, 'sp4_h_r_14')
// (19, 19, 'sp4_h_r_14')
// (20, 13, 'sp4_h_r_28')
// (20, 14, 'local_g2_0')
// (20, 14, 'local_g3_2')
// (20, 14, 'lutff_1/in_0')
// (20, 14, 'lutff_5/in_1')
// (20, 14, 'sp4_h_r_26')
// (20, 14, 'sp4_h_r_32')
// (20, 18, 'sp4_h_r_27')
// (20, 19, 'sp4_h_r_27')
// (21, 13, 'sp4_h_r_41')
// (21, 14, 'sp4_h_r_39')
// (21, 14, 'sp4_h_r_45')
// (21, 14, 'sp4_r_v_b_41')
// (21, 15, 'sp4_r_v_b_28')
// (21, 16, 'sp4_r_v_b_17')
// (21, 17, 'sp4_r_v_b_4')
// (21, 18, 'sp4_h_r_38')
// (21, 18, 'sp4_r_v_b_42')
// (21, 19, 'local_g1_7')
// (21, 19, 'local_g3_6')
// (21, 19, 'lutff_2/in_0')
// (21, 19, 'lutff_5/in_0')
// (21, 19, 'sp4_h_r_38')
// (21, 19, 'sp4_r_v_b_31')
// (21, 20, 'sp4_r_v_b_18')
// (21, 21, 'sp4_r_v_b_7')
// (22, 13, 'sp4_h_l_41')
// (22, 13, 'sp4_v_t_41')
// (22, 14, 'sp4_h_l_39')
// (22, 14, 'sp4_h_l_45')
// (22, 14, 'sp4_v_b_41')
// (22, 15, 'sp4_v_b_28')
// (22, 16, 'sp4_v_b_17')
// (22, 17, 'local_g0_4')
// (22, 17, 'lutff_0/in_2')
// (22, 17, 'lutff_6/in_2')
// (22, 17, 'sp4_v_b_4')
// (22, 17, 'sp4_v_t_42')
// (22, 18, 'local_g1_3')
// (22, 18, 'local_g1_6')
// (22, 18, 'lutff_1/in_0')
// (22, 18, 'lutff_6/in_0')
// (22, 18, 'sp4_h_l_38')
// (22, 18, 'sp4_h_r_3')
// (22, 18, 'sp4_h_r_6')
// (22, 18, 'sp4_v_b_42')
// (22, 19, 'sp4_h_l_38')
// (22, 19, 'sp4_v_b_31')
// (22, 20, 'sp4_v_b_18')
// (22, 21, 'sp4_v_b_7')
// (23, 18, 'sp4_h_r_14')
// (23, 18, 'sp4_h_r_19')
// (24, 18, 'sp4_h_r_27')
// (24, 18, 'sp4_h_r_30')
// (25, 18, 'sp4_h_r_38')
// (25, 18, 'sp4_h_r_43')
// (26, 18, 'sp4_h_l_38')
// (26, 18, 'sp4_h_l_43')

wire n706;
// (13, 16, 'neigh_op_tnr_0')
// (13, 17, 'local_g0_5')
// (13, 17, 'lutff_3/in_0')
// (13, 17, 'neigh_op_rgt_0')
// (13, 17, 'sp4_h_r_5')
// (13, 18, 'neigh_op_bnr_0')
// (14, 16, 'neigh_op_top_0')
// (14, 17, 'lutff_0/out')
// (14, 17, 'sp4_h_r_16')
// (14, 18, 'neigh_op_bot_0')
// (15, 16, 'neigh_op_tnl_0')
// (15, 17, 'neigh_op_lft_0')
// (15, 17, 'sp4_h_r_29')
// (15, 18, 'neigh_op_bnl_0')
// (16, 17, 'sp4_h_r_40')
// (17, 17, 'sp4_h_l_40')

wire n707;
// (13, 16, 'neigh_op_tnr_1')
// (13, 17, 'local_g3_1')
// (13, 17, 'lutff_3/in_1')
// (13, 17, 'neigh_op_rgt_1')
// (13, 18, 'neigh_op_bnr_1')
// (14, 16, 'neigh_op_top_1')
// (14, 17, 'lutff_1/out')
// (14, 18, 'neigh_op_bot_1')
// (15, 16, 'neigh_op_tnl_1')
// (15, 17, 'neigh_op_lft_1')
// (15, 18, 'neigh_op_bnl_1')

wire n708;
// (13, 16, 'neigh_op_tnr_2')
// (13, 17, 'local_g2_2')
// (13, 17, 'lutff_3/in_3')
// (13, 17, 'neigh_op_rgt_2')
// (13, 18, 'neigh_op_bnr_2')
// (14, 16, 'neigh_op_top_2')
// (14, 17, 'lutff_2/out')
// (14, 18, 'neigh_op_bot_2')
// (15, 16, 'neigh_op_tnl_2')
// (15, 17, 'neigh_op_lft_2')
// (15, 18, 'neigh_op_bnl_2')

reg n709 = 0;
// (13, 16, 'sp12_h_r_1')
// (14, 13, 'sp4_h_r_1')
// (14, 14, 'sp4_h_r_10')
// (14, 16, 'sp12_h_r_2')
// (15, 13, 'sp4_h_r_12')
// (15, 14, 'sp4_h_r_23')
// (15, 16, 'sp12_h_r_5')
// (16, 13, 'sp4_h_r_25')
// (16, 14, 'sp4_h_r_34')
// (16, 16, 'sp12_h_r_6')
// (17, 10, 'sp4_r_v_b_38')
// (17, 11, 'local_g0_3')
// (17, 11, 'lutff_2/in_1')
// (17, 11, 'lutff_4/in_1')
// (17, 11, 'sp4_r_v_b_27')
// (17, 12, 'sp4_r_v_b_14')
// (17, 13, 'local_g2_4')
// (17, 13, 'local_g3_4')
// (17, 13, 'lutff_3/in_2')
// (17, 13, 'lutff_4/in_0')
// (17, 13, 'sp4_h_r_36')
// (17, 13, 'sp4_r_v_b_3')
// (17, 14, 'sp4_h_r_47')
// (17, 14, 'sp4_r_v_b_42')
// (17, 15, 'neigh_op_tnr_1')
// (17, 15, 'sp4_r_v_b_31')
// (17, 15, 'sp4_r_v_b_47')
// (17, 16, 'local_g2_2')
// (17, 16, 'local_g3_2')
// (17, 16, 'lutff_5/in_1')
// (17, 16, 'lutff_6/in_1')
// (17, 16, 'neigh_op_rgt_1')
// (17, 16, 'sp12_h_r_9')
// (17, 16, 'sp4_r_v_b_18')
// (17, 16, 'sp4_r_v_b_34')
// (17, 17, 'local_g1_1')
// (17, 17, 'lutff_2/in_0')
// (17, 17, 'lutff_7/in_3')
// (17, 17, 'neigh_op_bnr_1')
// (17, 17, 'sp4_r_v_b_23')
// (17, 17, 'sp4_r_v_b_7')
// (17, 18, 'sp4_r_v_b_10')
// (17, 18, 'sp4_r_v_b_42')
// (17, 19, 'sp4_r_v_b_31')
// (17, 20, 'sp4_r_v_b_18')
// (17, 21, 'sp4_r_v_b_7')
// (18, 9, 'sp4_v_t_38')
// (18, 10, 'sp4_v_b_38')
// (18, 11, 'sp4_v_b_27')
// (18, 12, 'sp4_v_b_14')
// (18, 13, 'local_g0_3')
// (18, 13, 'local_g1_7')
// (18, 13, 'lutff_2/in_2')
// (18, 13, 'lutff_3/in_0')
// (18, 13, 'lutff_6/in_2')
// (18, 13, 'lutff_7/in_0')
// (18, 13, 'sp12_v_t_22')
// (18, 13, 'sp4_h_l_36')
// (18, 13, 'sp4_h_r_7')
// (18, 13, 'sp4_v_b_3')
// (18, 13, 'sp4_v_t_42')
// (18, 14, 'local_g2_2')
// (18, 14, 'local_g3_6')
// (18, 14, 'lutff_2/in_2')
// (18, 14, 'lutff_3/in_0')
// (18, 14, 'lutff_4/in_2')
// (18, 14, 'lutff_5/in_1')
// (18, 14, 'sp12_v_b_22')
// (18, 14, 'sp4_h_l_47')
// (18, 14, 'sp4_h_r_3')
// (18, 14, 'sp4_h_r_6')
// (18, 14, 'sp4_r_v_b_43')
// (18, 14, 'sp4_v_b_42')
// (18, 14, 'sp4_v_t_47')
// (18, 15, 'local_g3_7')
// (18, 15, 'lutff_6/in_0')
// (18, 15, 'neigh_op_top_1')
// (18, 15, 'sp12_v_b_21')
// (18, 15, 'sp4_r_v_b_30')
// (18, 15, 'sp4_v_b_31')
// (18, 15, 'sp4_v_b_47')
// (18, 16, 'local_g3_1')
// (18, 16, 'lutff_1/in_1')
// (18, 16, 'lutff_1/out')
// (18, 16, 'sp12_h_r_10')
// (18, 16, 'sp12_v_b_18')
// (18, 16, 'sp4_h_r_2')
// (18, 16, 'sp4_r_v_b_19')
// (18, 16, 'sp4_v_b_18')
// (18, 16, 'sp4_v_b_34')
// (18, 17, 'local_g0_1')
// (18, 17, 'local_g1_1')
// (18, 17, 'lutff_2/in_0')
// (18, 17, 'lutff_5/in_0')
// (18, 17, 'lutff_6/in_0')
// (18, 17, 'neigh_op_bot_1')
// (18, 17, 'sp12_v_b_17')
// (18, 17, 'sp4_h_r_7')
// (18, 17, 'sp4_r_v_b_6')
// (18, 17, 'sp4_v_b_23')
// (18, 17, 'sp4_v_b_7')
// (18, 17, 'sp4_v_t_42')
// (18, 18, 'local_g0_2')
// (18, 18, 'local_g3_2')
// (18, 18, 'lutff_2/in_0')
// (18, 18, 'lutff_6/in_0')
// (18, 18, 'lutff_7/in_0')
// (18, 18, 'sp12_v_b_14')
// (18, 18, 'sp4_h_r_4')
// (18, 18, 'sp4_r_v_b_43')
// (18, 18, 'sp4_v_b_10')
// (18, 18, 'sp4_v_b_42')
// (18, 19, 'sp12_v_b_13')
// (18, 19, 'sp4_r_v_b_30')
// (18, 19, 'sp4_v_b_31')
// (18, 20, 'local_g0_2')
// (18, 20, 'local_g1_2')
// (18, 20, 'lutff_1/in_1')
// (18, 20, 'lutff_2/in_0')
// (18, 20, 'lutff_7/in_2')
// (18, 20, 'sp12_v_b_10')
// (18, 20, 'sp4_r_v_b_19')
// (18, 20, 'sp4_v_b_18')
// (18, 21, 'sp12_v_b_9')
// (18, 21, 'sp4_h_r_7')
// (18, 21, 'sp4_r_v_b_6')
// (18, 21, 'sp4_v_b_7')
// (18, 22, 'sp12_v_b_6')
// (18, 23, 'sp12_v_b_5')
// (18, 24, 'local_g3_2')
// (18, 24, 'lutff_4/in_1')
// (18, 24, 'lutff_5/in_0')
// (18, 24, 'lutff_7/in_2')
// (18, 24, 'sp12_v_b_2')
// (18, 25, 'sp12_v_b_1')
// (19, 13, 'local_g1_2')
// (19, 13, 'lutff_3/in_0')
// (19, 13, 'sp4_h_r_18')
// (19, 13, 'sp4_v_t_43')
// (19, 14, 'local_g1_6')
// (19, 14, 'lutff_5/in_0')
// (19, 14, 'sp4_h_r_14')
// (19, 14, 'sp4_h_r_19')
// (19, 14, 'sp4_v_b_43')
// (19, 15, 'neigh_op_tnl_1')
// (19, 15, 'sp4_v_b_30')
// (19, 16, 'neigh_op_lft_1')
// (19, 16, 'sp12_h_r_13')
// (19, 16, 'sp4_h_r_15')
// (19, 16, 'sp4_v_b_19')
// (19, 17, 'local_g0_2')
// (19, 17, 'local_g2_1')
// (19, 17, 'lutff_0/in_2')
// (19, 17, 'lutff_3/in_2')
// (19, 17, 'lutff_4/in_2')
// (19, 17, 'lutff_5/in_0')
// (19, 17, 'neigh_op_bnl_1')
// (19, 17, 'sp4_h_r_18')
// (19, 17, 'sp4_v_b_6')
// (19, 17, 'sp4_v_t_43')
// (19, 18, 'local_g2_3')
// (19, 18, 'lutff_5/in_0')
// (19, 18, 'sp4_h_r_17')
// (19, 18, 'sp4_v_b_43')
// (19, 19, 'sp4_v_b_30')
// (19, 20, 'sp4_v_b_19')
// (19, 21, 'sp4_h_r_0')
// (19, 21, 'sp4_h_r_18')
// (19, 21, 'sp4_v_b_6')
// (20, 13, 'local_g3_7')
// (20, 13, 'lutff_2/in_0')
// (20, 13, 'lutff_4/in_0')
// (20, 13, 'sp4_h_r_31')
// (20, 14, 'local_g2_3')
// (20, 14, 'local_g2_6')
// (20, 14, 'lutff_0/in_2')
// (20, 14, 'lutff_3/in_2')
// (20, 14, 'lutff_4/in_0')
// (20, 14, 'lutff_6/in_2')
// (20, 14, 'sp4_h_r_27')
// (20, 14, 'sp4_h_r_30')
// (20, 16, 'sp12_h_r_14')
// (20, 16, 'sp4_h_r_26')
// (20, 17, 'sp4_h_r_31')
// (20, 18, 'sp4_h_r_28')
// (20, 21, 'sp4_h_r_13')
// (20, 21, 'sp4_h_r_31')
// (21, 13, 'local_g3_2')
// (21, 13, 'lutff_3/in_0')
// (21, 13, 'sp4_h_r_42')
// (21, 14, 'sp4_h_r_38')
// (21, 14, 'sp4_h_r_43')
// (21, 15, 'local_g3_1')
// (21, 15, 'lutff_2/in_0')
// (21, 15, 'lutff_4/in_0')
// (21, 15, 'sp4_r_v_b_41')
// (21, 16, 'local_g3_7')
// (21, 16, 'lutff_7/in_1')
// (21, 16, 'sp12_h_r_17')
// (21, 16, 'sp4_h_r_39')
// (21, 16, 'sp4_r_v_b_28')
// (21, 17, 'sp4_h_r_42')
// (21, 17, 'sp4_r_v_b_17')
// (21, 17, 'sp4_r_v_b_39')
// (21, 18, 'sp4_h_r_41')
// (21, 18, 'sp4_r_v_b_26')
// (21, 18, 'sp4_r_v_b_36')
// (21, 18, 'sp4_r_v_b_4')
// (21, 19, 'local_g2_7')
// (21, 19, 'local_g3_7')
// (21, 19, 'lutff_0/in_2')
// (21, 19, 'lutff_1/in_0')
// (21, 19, 'lutff_3/in_2')
// (21, 19, 'lutff_4/in_0')
// (21, 19, 'sp4_r_v_b_15')
// (21, 19, 'sp4_r_v_b_25')
// (21, 19, 'sp4_r_v_b_47')
// (21, 20, 'sp4_r_v_b_12')
// (21, 20, 'sp4_r_v_b_2')
// (21, 20, 'sp4_r_v_b_34')
// (21, 21, 'local_g2_2')
// (21, 21, 'local_g3_0')
// (21, 21, 'lutff_1/in_1')
// (21, 21, 'lutff_2/in_0')
// (21, 21, 'lutff_7/in_2')
// (21, 21, 'sp4_h_r_24')
// (21, 21, 'sp4_h_r_42')
// (21, 21, 'sp4_r_v_b_1')
// (21, 21, 'sp4_r_v_b_23')
// (21, 22, 'sp4_r_v_b_10')
// (22, 13, 'sp4_h_l_42')
// (22, 14, 'sp4_h_l_38')
// (22, 14, 'sp4_h_l_43')
// (22, 14, 'sp4_v_t_41')
// (22, 15, 'sp4_v_b_41')
// (22, 16, 'local_g1_2')
// (22, 16, 'lutff_7/in_0')
// (22, 16, 'sp12_h_r_18')
// (22, 16, 'sp4_h_l_39')
// (22, 16, 'sp4_v_b_28')
// (22, 16, 'sp4_v_t_39')
// (22, 17, 'local_g0_1')
// (22, 17, 'local_g1_1')
// (22, 17, 'lutff_2/in_2')
// (22, 17, 'lutff_3/in_0')
// (22, 17, 'lutff_4/in_2')
// (22, 17, 'lutff_5/in_0')
// (22, 17, 'sp4_h_l_42')
// (22, 17, 'sp4_v_b_17')
// (22, 17, 'sp4_v_b_39')
// (22, 17, 'sp4_v_t_36')
// (22, 18, 'local_g2_4')
// (22, 18, 'local_g3_4')
// (22, 18, 'lutff_0/in_2')
// (22, 18, 'lutff_3/in_2')
// (22, 18, 'lutff_4/in_2')
// (22, 18, 'lutff_5/in_0')
// (22, 18, 'sp4_h_l_41')
// (22, 18, 'sp4_h_r_4')
// (22, 18, 'sp4_v_b_26')
// (22, 18, 'sp4_v_b_36')
// (22, 18, 'sp4_v_b_4')
// (22, 18, 'sp4_v_t_47')
// (22, 19, 'sp4_v_b_15')
// (22, 19, 'sp4_v_b_25')
// (22, 19, 'sp4_v_b_47')
// (22, 20, 'local_g0_4')
// (22, 20, 'local_g1_4')
// (22, 20, 'lutff_0/in_2')
// (22, 20, 'lutff_3/in_0')
// (22, 20, 'lutff_4/in_1')
// (22, 20, 'sp4_v_b_12')
// (22, 20, 'sp4_v_b_2')
// (22, 20, 'sp4_v_b_34')
// (22, 21, 'sp4_h_l_42')
// (22, 21, 'sp4_h_r_37')
// (22, 21, 'sp4_v_b_1')
// (22, 21, 'sp4_v_b_23')
// (22, 22, 'sp4_v_b_10')
// (23, 16, 'sp12_h_r_21')
// (23, 18, 'sp4_h_r_17')
// (23, 21, 'sp4_h_l_37')
// (24, 16, 'sp12_h_r_22')
// (24, 18, 'sp4_h_r_28')
// (25, 16, 'sp12_h_l_22')
// (25, 18, 'sp4_h_r_41')
// (26, 18, 'sp4_h_l_41')

wire n710;
// (13, 17, 'lutff_2/lout')
// (13, 17, 'lutff_3/in_2')

wire n711;
// (13, 17, 'lutff_3/lout')
// (13, 17, 'lutff_4/in_2')

wire n712;
// (13, 17, 'sp4_h_r_0')
// (14, 17, 'local_g1_5')
// (14, 17, 'lutff_5/in_3')
// (14, 17, 'sp4_h_r_13')
// (15, 17, 'sp4_h_r_24')
// (16, 14, 'sp4_r_v_b_41')
// (16, 15, 'sp4_r_v_b_28')
// (16, 16, 'sp4_r_v_b_17')
// (16, 17, 'sp4_h_r_37')
// (16, 17, 'sp4_r_v_b_4')
// (16, 18, 'sp4_r_v_b_37')
// (16, 18, 'sp4_r_v_b_45')
// (16, 19, 'sp4_r_v_b_24')
// (16, 19, 'sp4_r_v_b_32')
// (16, 20, 'sp4_r_v_b_13')
// (16, 20, 'sp4_r_v_b_21')
// (16, 21, 'sp4_r_v_b_0')
// (16, 21, 'sp4_r_v_b_8')
// (16, 22, 'sp4_r_v_b_37')
// (16, 23, 'sp4_r_v_b_24')
// (16, 24, 'neigh_op_tnr_0')
// (16, 24, 'sp4_r_v_b_13')
// (16, 25, 'neigh_op_rgt_0')
// (16, 25, 'sp4_r_v_b_0')
// (16, 26, 'neigh_op_bnr_0')
// (17, 9, 'sp12_v_t_23')
// (17, 10, 'local_g2_7')
// (17, 10, 'lutff_0/in_3')
// (17, 10, 'sp12_v_b_23')
// (17, 11, 'sp12_v_b_20')
// (17, 12, 'sp12_v_b_19')
// (17, 13, 'sp12_v_b_16')
// (17, 13, 'sp4_h_r_4')
// (17, 13, 'sp4_v_t_41')
// (17, 14, 'sp12_v_b_15')
// (17, 14, 'sp4_v_b_41')
// (17, 15, 'sp12_v_b_12')
// (17, 15, 'sp4_r_v_b_41')
// (17, 15, 'sp4_r_v_b_42')
// (17, 15, 'sp4_v_b_28')
// (17, 16, 'sp12_v_b_11')
// (17, 16, 'sp4_r_v_b_28')
// (17, 16, 'sp4_r_v_b_31')
// (17, 16, 'sp4_v_b_17')
// (17, 17, 'sp12_v_b_8')
// (17, 17, 'sp4_h_l_37')
// (17, 17, 'sp4_h_r_0')
// (17, 17, 'sp4_r_v_b_17')
// (17, 17, 'sp4_r_v_b_18')
// (17, 17, 'sp4_v_b_4')
// (17, 17, 'sp4_v_t_37')
// (17, 17, 'sp4_v_t_45')
// (17, 18, 'sp12_v_b_7')
// (17, 18, 'sp4_r_v_b_4')
// (17, 18, 'sp4_r_v_b_7')
// (17, 18, 'sp4_v_b_37')
// (17, 18, 'sp4_v_b_45')
// (17, 19, 'sp12_v_b_4')
// (17, 19, 'sp4_r_v_b_41')
// (17, 19, 'sp4_v_b_24')
// (17, 19, 'sp4_v_b_32')
// (17, 20, 'sp12_v_b_3')
// (17, 20, 'sp4_r_v_b_28')
// (17, 20, 'sp4_v_b_13')
// (17, 20, 'sp4_v_b_21')
// (17, 21, 'sp12_v_b_0')
// (17, 21, 'sp12_v_t_23')
// (17, 21, 'sp4_r_v_b_17')
// (17, 21, 'sp4_v_b_0')
// (17, 21, 'sp4_v_b_8')
// (17, 21, 'sp4_v_t_37')
// (17, 22, 'sp12_v_b_23')
// (17, 22, 'sp4_r_v_b_36')
// (17, 22, 'sp4_r_v_b_4')
// (17, 22, 'sp4_v_b_37')
// (17, 23, 'sp12_v_b_20')
// (17, 23, 'sp4_r_v_b_25')
// (17, 23, 'sp4_r_v_b_41')
// (17, 23, 'sp4_v_b_24')
// (17, 24, 'neigh_op_top_0')
// (17, 24, 'sp12_v_b_19')
// (17, 24, 'sp4_r_v_b_12')
// (17, 24, 'sp4_r_v_b_28')
// (17, 24, 'sp4_v_b_13')
// (17, 25, 'local_g0_0')
// (17, 25, 'lutff_0/out')
// (17, 25, 'lutff_1/in_1')
// (17, 25, 'sp12_v_b_16')
// (17, 25, 'sp4_r_v_b_1')
// (17, 25, 'sp4_r_v_b_17')
// (17, 25, 'sp4_v_b_0')
// (17, 26, 'neigh_op_bot_0')
// (17, 26, 'sp12_v_b_15')
// (17, 26, 'sp4_r_v_b_4')
// (17, 27, 'sp12_v_b_12')
// (17, 28, 'sp12_v_b_11')
// (17, 29, 'sp12_v_b_8')
// (17, 30, 'sp12_v_b_7')
// (17, 31, 'sp12_v_b_4')
// (17, 32, 'sp12_v_b_3')
// (17, 33, 'span12_vert_0')
// (18, 13, 'local_g1_1')
// (18, 13, 'lutff_1/in_3')
// (18, 13, 'sp4_h_r_17')
// (18, 14, 'local_g1_0')
// (18, 14, 'lutff_6/in_3')
// (18, 14, 'sp4_h_r_0')
// (18, 14, 'sp4_v_t_41')
// (18, 14, 'sp4_v_t_42')
// (18, 15, 'sp4_v_b_41')
// (18, 15, 'sp4_v_b_42')
// (18, 16, 'local_g3_4')
// (18, 16, 'local_g3_7')
// (18, 16, 'lutff_1/in_0')
// (18, 16, 'lutff_2/in_0')
// (18, 16, 'lutff_3/in_0')
// (18, 16, 'lutff_4/in_1')
// (18, 16, 'sp4_v_b_28')
// (18, 16, 'sp4_v_b_31')
// (18, 17, 'sp4_h_r_13')
// (18, 17, 'sp4_v_b_17')
// (18, 17, 'sp4_v_b_18')
// (18, 18, 'sp4_v_b_4')
// (18, 18, 'sp4_v_b_7')
// (18, 18, 'sp4_v_t_41')
// (18, 19, 'sp4_v_b_41')
// (18, 20, 'sp4_v_b_28')
// (18, 21, 'sp4_h_r_6')
// (18, 21, 'sp4_v_b_17')
// (18, 21, 'sp4_v_t_36')
// (18, 22, 'sp4_h_r_9')
// (18, 22, 'sp4_v_b_36')
// (18, 22, 'sp4_v_b_4')
// (18, 22, 'sp4_v_t_41')
// (18, 23, 'sp4_v_b_25')
// (18, 23, 'sp4_v_b_41')
// (18, 24, 'neigh_op_tnl_0')
// (18, 24, 'sp4_v_b_12')
// (18, 24, 'sp4_v_b_28')
// (18, 25, 'neigh_op_lft_0')
// (18, 25, 'sp4_v_b_1')
// (18, 25, 'sp4_v_b_17')
// (18, 26, 'neigh_op_bnl_0')
// (18, 26, 'sp4_v_b_4')
// (19, 13, 'sp4_h_r_28')
// (19, 14, 'sp4_h_r_13')
// (19, 17, 'local_g3_0')
// (19, 17, 'lutff_2/in_3')
// (19, 17, 'sp4_h_r_24')
// (19, 21, 'sp4_h_r_19')
// (19, 22, 'sp4_h_r_20')
// (20, 13, 'sp4_h_r_41')
// (20, 14, 'local_g3_0')
// (20, 14, 'lutff_2/in_3')
// (20, 14, 'sp4_h_r_24')
// (20, 17, 'sp4_h_r_37')
// (20, 21, 'sp4_h_r_30')
// (20, 22, 'sp4_h_r_33')
// (21, 13, 'sp4_h_l_41')
// (21, 14, 'sp4_h_r_37')
// (21, 17, 'sp4_h_l_37')
// (21, 17, 'sp4_h_r_0')
// (21, 18, 'sp4_r_v_b_43')
// (21, 19, 'local_g3_4')
// (21, 19, 'lutff_6/in_3')
// (21, 19, 'sp4_r_v_b_30')
// (21, 19, 'sp4_r_v_b_44')
// (21, 20, 'sp4_r_v_b_19')
// (21, 20, 'sp4_r_v_b_33')
// (21, 21, 'sp4_h_r_43')
// (21, 21, 'sp4_r_v_b_20')
// (21, 21, 'sp4_r_v_b_6')
// (21, 22, 'sp4_h_r_44')
// (21, 22, 'sp4_r_v_b_9')
// (22, 14, 'sp4_h_l_37')
// (22, 17, 'local_g1_5')
// (22, 17, 'lutff_1/in_3')
// (22, 17, 'sp4_h_r_13')
// (22, 17, 'sp4_v_t_43')
// (22, 18, 'local_g2_3')
// (22, 18, 'lutff_2/in_3')
// (22, 18, 'sp4_v_b_43')
// (22, 18, 'sp4_v_t_44')
// (22, 19, 'sp4_v_b_30')
// (22, 19, 'sp4_v_b_44')
// (22, 20, 'sp4_v_b_19')
// (22, 20, 'sp4_v_b_33')
// (22, 21, 'sp4_h_l_43')
// (22, 21, 'sp4_v_b_20')
// (22, 21, 'sp4_v_b_6')
// (22, 22, 'sp4_h_l_44')
// (22, 22, 'sp4_v_b_9')
// (23, 17, 'sp4_h_r_24')
// (24, 17, 'sp4_h_r_37')
// (25, 17, 'sp4_h_l_37')

wire n713;
// (13, 17, 'sp4_h_r_1')
// (14, 17, 'local_g1_4')
// (14, 17, 'lutff_4/in_3')
// (14, 17, 'sp4_h_r_12')
// (15, 17, 'sp4_h_r_25')
// (16, 14, 'sp4_r_v_b_36')
// (16, 15, 'neigh_op_tnr_6')
// (16, 15, 'sp4_r_v_b_25')
// (16, 16, 'neigh_op_rgt_6')
// (16, 16, 'sp4_r_v_b_12')
// (16, 17, 'neigh_op_bnr_6')
// (16, 17, 'sp4_h_r_36')
// (16, 17, 'sp4_r_v_b_1')
// (17, 13, 'sp4_v_t_36')
// (17, 14, 'sp4_v_b_36')
// (17, 15, 'neigh_op_top_6')
// (17, 15, 'sp4_v_b_25')
// (17, 16, 'lutff_6/out')
// (17, 16, 'sp4_v_b_12')
// (17, 17, 'neigh_op_bot_6')
// (17, 17, 'sp4_h_l_36')
// (17, 17, 'sp4_v_b_1')
// (18, 15, 'neigh_op_tnl_6')
// (18, 16, 'neigh_op_lft_6')
// (18, 17, 'neigh_op_bnl_6')

reg n714 = 0;
// (13, 17, 'sp4_h_r_2')
// (14, 16, 'neigh_op_tnr_5')
// (14, 17, 'neigh_op_rgt_5')
// (14, 17, 'sp4_h_r_15')
// (14, 18, 'neigh_op_bnr_5')
// (15, 16, 'neigh_op_top_5')
// (15, 17, 'lutff_5/out')
// (15, 17, 'sp4_h_r_26')
// (15, 18, 'neigh_op_bot_5')
// (16, 14, 'sp4_r_v_b_45')
// (16, 15, 'sp4_r_v_b_32')
// (16, 16, 'neigh_op_tnl_5')
// (16, 16, 'sp4_r_v_b_21')
// (16, 17, 'neigh_op_lft_5')
// (16, 17, 'sp4_h_r_39')
// (16, 17, 'sp4_r_v_b_8')
// (16, 18, 'neigh_op_bnl_5')
// (17, 13, 'sp4_v_t_45')
// (17, 14, 'local_g2_5')
// (17, 14, 'lutff_1/in_0')
// (17, 14, 'sp4_v_b_45')
// (17, 15, 'sp4_v_b_32')
// (17, 16, 'sp4_v_b_21')
// (17, 17, 'sp4_h_l_39')
// (17, 17, 'sp4_v_b_8')

wire n715;
// (13, 18, 'lutff_7/cout')
// (13, 19, 'carry_in')
// (13, 19, 'carry_in_mux')

reg n716 = 0;
// (13, 18, 'sp4_h_r_10')
// (14, 17, 'neigh_op_tnr_1')
// (14, 18, 'neigh_op_rgt_1')
// (14, 18, 'sp4_h_r_23')
// (14, 19, 'neigh_op_bnr_1')
// (15, 17, 'neigh_op_top_1')
// (15, 18, 'lutff_1/out')
// (15, 18, 'sp4_h_r_34')
// (15, 19, 'neigh_op_bot_1')
// (16, 17, 'neigh_op_tnl_1')
// (16, 18, 'neigh_op_lft_1')
// (16, 18, 'sp4_h_r_47')
// (16, 19, 'neigh_op_bnl_1')
// (17, 18, 'sp4_h_l_47')
// (17, 18, 'sp4_h_r_1')
// (18, 18, 'sp4_h_r_12')
// (19, 18, 'sp4_h_r_25')
// (20, 18, 'sp4_h_r_36')
// (20, 19, 'sp4_r_v_b_36')
// (20, 20, 'sp4_r_v_b_25')
// (20, 21, 'sp4_r_v_b_12')
// (20, 22, 'sp4_r_v_b_1')
// (21, 18, 'sp4_h_l_36')
// (21, 18, 'sp4_v_t_36')
// (21, 19, 'sp4_v_b_36')
// (21, 20, 'sp4_v_b_25')
// (21, 21, 'local_g0_4')
// (21, 21, 'lutff_5/in_1')
// (21, 21, 'sp4_v_b_12')
// (21, 22, 'sp4_v_b_1')

wire n717;
// (13, 19, 'lutff_7/cout')
// (13, 20, 'carry_in')
// (13, 20, 'carry_in_mux')

reg n718 = 0;
// (13, 19, 'sp4_r_v_b_45')
// (13, 20, 'sp4_r_v_b_32')
// (13, 21, 'neigh_op_tnr_4')
// (13, 21, 'sp4_r_v_b_21')
// (13, 22, 'neigh_op_rgt_4')
// (13, 22, 'sp4_r_v_b_8')
// (13, 23, 'neigh_op_bnr_4')
// (14, 18, 'sp4_h_r_8')
// (14, 18, 'sp4_v_t_45')
// (14, 19, 'sp4_v_b_45')
// (14, 20, 'sp4_v_b_32')
// (14, 21, 'neigh_op_top_4')
// (14, 21, 'sp4_v_b_21')
// (14, 22, 'lutff_4/out')
// (14, 22, 'sp4_v_b_8')
// (14, 23, 'neigh_op_bot_4')
// (15, 18, 'sp4_h_r_21')
// (15, 21, 'neigh_op_tnl_4')
// (15, 22, 'neigh_op_lft_4')
// (15, 23, 'neigh_op_bnl_4')
// (16, 18, 'sp4_h_r_32')
// (17, 18, 'sp4_h_r_45')
// (18, 18, 'local_g1_3')
// (18, 18, 'lutff_5/in_3')
// (18, 18, 'sp4_h_l_45')
// (18, 18, 'sp4_h_r_11')
// (19, 18, 'sp4_h_r_22')
// (20, 18, 'sp4_h_r_35')
// (21, 18, 'sp4_h_r_46')
// (22, 18, 'sp4_h_l_46')

wire n719;
// (13, 20, 'lutff_7/cout')
// (13, 21, 'carry_in')
// (13, 21, 'carry_in_mux')
// (13, 21, 'lutff_0/in_3')

reg n720 = 0;
// (13, 20, 'neigh_op_tnr_6')
// (13, 21, 'neigh_op_rgt_6')
// (13, 22, 'neigh_op_bnr_6')
// (14, 20, 'neigh_op_top_6')
// (14, 21, 'lutff_6/out')
// (14, 22, 'neigh_op_bot_6')
// (15, 20, 'local_g3_6')
// (15, 20, 'lutff_2/in_3')
// (15, 20, 'neigh_op_tnl_6')
// (15, 21, 'neigh_op_lft_6')
// (15, 22, 'neigh_op_bnl_6')

reg n721 = 0;
// (13, 20, 'sp12_h_r_1')
// (14, 20, 'sp12_h_r_2')
// (15, 20, 'sp12_h_r_5')
// (16, 20, 'sp12_h_r_6')
// (17, 20, 'sp12_h_r_9')
// (18, 20, 'sp12_h_r_10')
// (19, 19, 'neigh_op_tnr_3')
// (19, 20, 'neigh_op_rgt_3')
// (19, 20, 'sp12_h_r_13')
// (19, 21, 'neigh_op_bnr_3')
// (20, 19, 'neigh_op_top_3')
// (20, 20, 'lutff_3/out')
// (20, 20, 'sp12_h_r_14')
// (20, 21, 'neigh_op_bot_3')
// (21, 19, 'neigh_op_tnl_3')
// (21, 20, 'neigh_op_lft_3')
// (21, 20, 'sp12_h_r_17')
// (21, 21, 'neigh_op_bnl_3')
// (22, 20, 'local_g1_2')
// (22, 20, 'lutff_2/in_1')
// (22, 20, 'sp12_h_r_18')
// (23, 20, 'sp12_h_r_21')
// (24, 20, 'sp12_h_r_22')
// (25, 20, 'sp12_h_l_22')

reg n722 = 0;
// (13, 21, 'neigh_op_tnr_0')
// (13, 21, 'sp4_r_v_b_45')
// (13, 22, 'neigh_op_rgt_0')
// (13, 22, 'sp4_r_v_b_32')
// (13, 23, 'neigh_op_bnr_0')
// (13, 23, 'sp4_r_v_b_21')
// (13, 24, 'sp4_r_v_b_8')
// (14, 20, 'sp4_h_r_1')
// (14, 20, 'sp4_v_t_45')
// (14, 21, 'neigh_op_top_0')
// (14, 21, 'sp4_v_b_45')
// (14, 22, 'lutff_0/out')
// (14, 22, 'sp4_v_b_32')
// (14, 23, 'neigh_op_bot_0')
// (14, 23, 'sp4_v_b_21')
// (14, 24, 'sp4_v_b_8')
// (15, 20, 'sp4_h_r_12')
// (15, 21, 'neigh_op_tnl_0')
// (15, 22, 'neigh_op_lft_0')
// (15, 23, 'neigh_op_bnl_0')
// (16, 20, 'sp4_h_r_25')
// (17, 17, 'sp4_r_v_b_42')
// (17, 18, 'sp4_r_v_b_31')
// (17, 19, 'sp4_r_v_b_18')
// (17, 20, 'sp4_h_r_36')
// (17, 20, 'sp4_r_v_b_7')
// (18, 16, 'sp4_v_t_42')
// (18, 17, 'local_g3_2')
// (18, 17, 'lutff_4/in_3')
// (18, 17, 'sp4_v_b_42')
// (18, 18, 'sp4_v_b_31')
// (18, 19, 'sp4_v_b_18')
// (18, 20, 'sp4_h_l_36')
// (18, 20, 'sp4_v_b_7')

reg n723 = 0;
// (13, 21, 'neigh_op_tnr_2')
// (13, 22, 'neigh_op_rgt_2')
// (13, 23, 'neigh_op_bnr_2')
// (14, 20, 'sp12_h_r_0')
// (14, 20, 'sp12_v_t_23')
// (14, 21, 'neigh_op_top_2')
// (14, 21, 'sp12_v_b_23')
// (14, 22, 'lutff_2/out')
// (14, 22, 'sp12_v_b_20')
// (14, 23, 'neigh_op_bot_2')
// (14, 23, 'sp12_v_b_19')
// (14, 24, 'sp12_v_b_16')
// (14, 25, 'sp12_v_b_15')
// (14, 26, 'sp12_v_b_12')
// (14, 27, 'sp12_v_b_11')
// (14, 28, 'sp12_v_b_8')
// (14, 29, 'sp12_v_b_7')
// (14, 30, 'sp12_v_b_4')
// (14, 31, 'sp12_v_b_3')
// (14, 32, 'sp12_v_b_0')
// (15, 20, 'sp12_h_r_3')
// (15, 21, 'neigh_op_tnl_2')
// (15, 22, 'neigh_op_lft_2')
// (15, 23, 'neigh_op_bnl_2')
// (16, 20, 'sp12_h_r_4')
// (17, 20, 'sp12_h_r_7')
// (18, 20, 'sp12_h_r_8')
// (19, 20, 'sp12_h_r_11')
// (20, 20, 'sp12_h_r_12')
// (21, 20, 'sp12_h_r_15')
// (22, 20, 'local_g1_0')
// (22, 20, 'lutff_2/in_3')
// (22, 20, 'sp12_h_r_16')
// (23, 20, 'sp12_h_r_19')
// (24, 20, 'sp12_h_r_20')
// (25, 20, 'sp12_h_r_23')
// (26, 20, 'sp12_h_l_23')

reg n724 = 0;
// (13, 21, 'neigh_op_tnr_3')
// (13, 22, 'neigh_op_rgt_3')
// (13, 22, 'sp4_r_v_b_38')
// (13, 23, 'neigh_op_bnr_3')
// (13, 23, 'sp4_r_v_b_27')
// (13, 24, 'sp4_r_v_b_14')
// (13, 25, 'sp4_r_v_b_3')
// (14, 21, 'neigh_op_top_3')
// (14, 21, 'sp4_h_r_3')
// (14, 21, 'sp4_v_t_38')
// (14, 22, 'lutff_3/out')
// (14, 22, 'sp4_v_b_38')
// (14, 23, 'neigh_op_bot_3')
// (14, 23, 'sp4_v_b_27')
// (14, 24, 'sp4_v_b_14')
// (14, 25, 'sp4_v_b_3')
// (15, 21, 'neigh_op_tnl_3')
// (15, 21, 'sp4_h_r_14')
// (15, 22, 'neigh_op_lft_3')
// (15, 23, 'neigh_op_bnl_3')
// (16, 21, 'sp4_h_r_27')
// (17, 21, 'local_g2_6')
// (17, 21, 'lutff_5/in_3')
// (17, 21, 'sp4_h_r_38')
// (18, 21, 'sp4_h_l_38')

reg n725 = 0;
// (13, 21, 'neigh_op_tnr_5')
// (13, 22, 'neigh_op_rgt_5')
// (13, 23, 'neigh_op_bnr_5')
// (14, 21, 'neigh_op_top_5')
// (14, 22, 'lutff_5/out')
// (14, 22, 'sp4_r_v_b_43')
// (14, 23, 'neigh_op_bot_5')
// (14, 23, 'sp4_r_v_b_30')
// (14, 24, 'sp4_r_v_b_19')
// (14, 25, 'sp4_r_v_b_6')
// (15, 21, 'neigh_op_tnl_5')
// (15, 21, 'sp4_v_t_43')
// (15, 22, 'neigh_op_lft_5')
// (15, 22, 'sp4_v_b_43')
// (15, 23, 'neigh_op_bnl_5')
// (15, 23, 'sp4_v_b_30')
// (15, 24, 'sp4_v_b_19')
// (15, 25, 'sp4_h_r_6')
// (15, 25, 'sp4_v_b_6')
// (16, 25, 'sp4_h_r_19')
// (17, 25, 'sp4_h_r_30')
// (18, 25, 'local_g3_3')
// (18, 25, 'lutff_5/in_3')
// (18, 25, 'sp4_h_r_43')
// (19, 25, 'sp4_h_l_43')

reg io_33_23_1 = 0;
// (13, 21, 'sp12_h_r_1')
// (14, 21, 'sp12_h_r_2')
// (15, 21, 'sp12_h_r_5')
// (16, 21, 'sp12_h_r_6')
// (17, 20, 'neigh_op_tnr_1')
// (17, 21, 'neigh_op_rgt_1')
// (17, 21, 'sp12_h_r_9')
// (17, 22, 'neigh_op_bnr_1')
// (18, 20, 'neigh_op_top_1')
// (18, 21, 'lutff_1/out')
// (18, 21, 'sp12_h_r_10')
// (18, 22, 'neigh_op_bot_1')
// (19, 20, 'neigh_op_tnl_1')
// (19, 21, 'neigh_op_lft_1')
// (19, 21, 'sp12_h_r_13')
// (19, 22, 'neigh_op_bnl_1')
// (20, 21, 'sp12_h_r_14')
// (21, 21, 'sp12_h_r_17')
// (22, 21, 'sp12_h_r_18')
// (23, 21, 'sp12_h_r_21')
// (24, 21, 'sp12_h_r_22')
// (25, 21, 'sp12_h_l_22')
// (25, 21, 'sp12_h_r_1')
// (26, 21, 'sp12_h_r_2')
// (27, 21, 'sp12_h_r_5')
// (28, 21, 'sp12_h_r_6')
// (29, 21, 'sp12_h_r_9')
// (30, 21, 'sp12_h_r_10')
// (31, 21, 'sp12_h_r_13')
// (31, 21, 'sp4_h_r_6')
// (32, 21, 'sp12_h_r_14')
// (32, 21, 'sp4_h_r_19')
// (33, 21, 'span12_horz_14')
// (33, 21, 'span4_horz_19')
// (33, 21, 'span4_vert_t_15')
// (33, 22, 'span4_vert_b_15')
// (33, 23, 'io_1/D_OUT_0')
// (33, 23, 'io_1/PAD')
// (33, 23, 'local_g0_3')
// (33, 23, 'span4_vert_b_11')
// (33, 24, 'span4_vert_b_7')
// (33, 25, 'span4_vert_b_3')

wire n727;
// (13, 22, 'lutff_7/cout')
// (13, 23, 'carry_in')
// (13, 23, 'carry_in_mux')

wire n728;
// (13, 23, 'lutff_7/cout')
// (13, 24, 'carry_in')
// (13, 24, 'carry_in_mux')

reg n729 = 0;
// (13, 23, 'sp12_h_r_0')
// (14, 23, 'sp12_h_r_3')
// (15, 23, 'sp12_h_r_4')
// (16, 23, 'sp12_h_r_7')
// (17, 23, 'sp12_h_r_8')
// (18, 22, 'neigh_op_tnr_2')
// (18, 23, 'neigh_op_rgt_2')
// (18, 23, 'sp12_h_r_11')
// (18, 24, 'neigh_op_bnr_2')
// (19, 22, 'neigh_op_top_2')
// (19, 23, 'local_g2_2')
// (19, 23, 'lutff_2/in_0')
// (19, 23, 'lutff_2/out')
// (19, 23, 'sp12_h_r_12')
// (19, 24, 'neigh_op_bot_2')
// (20, 22, 'neigh_op_tnl_2')
// (20, 23, 'neigh_op_lft_2')
// (20, 23, 'sp12_h_r_15')
// (20, 24, 'neigh_op_bnl_2')
// (21, 23, 'sp12_h_r_16')
// (22, 23, 'sp12_h_r_19')
// (23, 23, 'sp12_h_r_20')
// (24, 23, 'sp12_h_r_23')
// (25, 23, 'sp12_h_l_23')
// (25, 23, 'sp12_h_r_0')
// (26, 23, 'sp12_h_r_3')
// (27, 23, 'sp12_h_r_4')
// (28, 23, 'sp12_h_r_7')
// (29, 23, 'sp12_h_r_8')
// (30, 23, 'sp12_h_r_11')
// (30, 23, 'sp4_h_r_7')
// (31, 23, 'sp12_h_r_12')
// (31, 23, 'sp4_h_r_18')
// (32, 23, 'sp12_h_r_15')
// (32, 23, 'sp4_h_r_31')
// (33, 15, 'span4_vert_t_13')
// (33, 16, 'io_1/OUT_ENB')
// (33, 16, 'local_g1_5')
// (33, 16, 'span4_vert_b_13')
// (33, 17, 'span4_vert_b_9')
// (33, 18, 'span4_vert_b_5')
// (33, 19, 'span4_vert_b_1')
// (33, 19, 'span4_vert_t_13')
// (33, 20, 'span4_vert_b_13')
// (33, 21, 'span4_vert_b_9')
// (33, 22, 'span4_vert_b_5')
// (33, 23, 'span12_horz_15')
// (33, 23, 'span4_horz_31')
// (33, 23, 'span4_vert_b_1')

reg io_33_29_1 = 0;
// (13, 23, 'sp12_h_r_1')
// (14, 23, 'sp12_h_r_2')
// (15, 23, 'sp12_h_r_5')
// (16, 23, 'sp12_h_r_6')
// (17, 22, 'neigh_op_tnr_1')
// (17, 23, 'neigh_op_rgt_1')
// (17, 23, 'sp12_h_r_9')
// (17, 24, 'neigh_op_bnr_1')
// (18, 22, 'neigh_op_top_1')
// (18, 23, 'lutff_1/out')
// (18, 23, 'sp12_h_r_10')
// (18, 24, 'neigh_op_bot_1')
// (19, 22, 'neigh_op_tnl_1')
// (19, 23, 'neigh_op_lft_1')
// (19, 23, 'sp12_h_r_13')
// (19, 24, 'neigh_op_bnl_1')
// (20, 23, 'sp12_h_r_14')
// (21, 23, 'sp12_h_r_17')
// (22, 23, 'sp12_h_r_18')
// (23, 23, 'sp12_h_r_21')
// (24, 23, 'sp12_h_r_22')
// (25, 23, 'sp12_h_l_22')
// (25, 23, 'sp12_h_r_1')
// (26, 23, 'sp12_h_r_2')
// (27, 23, 'sp12_h_r_5')
// (28, 23, 'sp12_h_r_6')
// (29, 23, 'sp12_h_r_9')
// (30, 23, 'sp12_h_r_10')
// (31, 23, 'sp12_h_r_13')
// (31, 23, 'sp4_h_r_6')
// (32, 23, 'sp12_h_r_14')
// (32, 23, 'sp4_h_r_19')
// (33, 23, 'span12_horz_14')
// (33, 23, 'span4_horz_19')
// (33, 23, 'span4_vert_t_15')
// (33, 24, 'span4_vert_b_15')
// (33, 25, 'span4_vert_b_11')
// (33, 26, 'span4_vert_b_7')
// (33, 27, 'span4_vert_b_3')
// (33, 27, 'span4_vert_t_15')
// (33, 28, 'span4_vert_b_15')
// (33, 29, 'io_1/D_OUT_0')
// (33, 29, 'io_1/PAD')
// (33, 29, 'local_g0_3')
// (33, 29, 'span4_vert_b_11')
// (33, 30, 'span4_vert_b_7')
// (33, 31, 'span4_vert_b_3')

wire n731;
// (13, 23, 'sp4_h_r_8')
// (14, 22, 'neigh_op_tnr_0')
// (14, 23, 'neigh_op_rgt_0')
// (14, 23, 'sp4_h_r_21')
// (14, 23, 'sp4_h_r_5')
// (14, 24, 'neigh_op_bnr_0')
// (15, 22, 'neigh_op_top_0')
// (15, 22, 'sp4_r_v_b_44')
// (15, 23, 'lutff_0/out')
// (15, 23, 'sp4_h_r_16')
// (15, 23, 'sp4_h_r_32')
// (15, 23, 'sp4_r_v_b_33')
// (15, 24, 'neigh_op_bot_0')
// (15, 24, 'sp4_r_v_b_20')
// (15, 25, 'sp4_r_v_b_9')
// (16, 21, 'sp4_h_r_9')
// (16, 21, 'sp4_v_t_44')
// (16, 22, 'local_g2_0')
// (16, 22, 'lutff_0/in_0')
// (16, 22, 'lutff_1/in_3')
// (16, 22, 'lutff_2/in_0')
// (16, 22, 'lutff_3/in_3')
// (16, 22, 'lutff_4/in_0')
// (16, 22, 'neigh_op_tnl_0')
// (16, 22, 'sp4_v_b_44')
// (16, 23, 'neigh_op_lft_0')
// (16, 23, 'sp4_h_r_29')
// (16, 23, 'sp4_h_r_45')
// (16, 23, 'sp4_v_b_33')
// (16, 24, 'neigh_op_bnl_0')
// (16, 24, 'sp4_v_b_20')
// (16, 25, 'sp4_v_b_9')
// (17, 20, 'sp4_r_v_b_40')
// (17, 21, 'sp4_h_r_20')
// (17, 21, 'sp4_r_v_b_29')
// (17, 22, 'sp4_r_v_b_16')
// (17, 23, 'sp4_h_l_45')
// (17, 23, 'sp4_h_r_40')
// (17, 23, 'sp4_h_r_8')
// (17, 23, 'sp4_r_v_b_5')
// (18, 19, 'sp4_v_t_40')
// (18, 20, 'sp4_v_b_40')
// (18, 21, 'local_g2_5')
// (18, 21, 'local_g3_1')
// (18, 21, 'lutff_0/in_3')
// (18, 21, 'lutff_1/in_0')
// (18, 21, 'lutff_2/in_1')
// (18, 21, 'lutff_3/in_1')
// (18, 21, 'lutff_4/in_3')
// (18, 21, 'lutff_5/in_0')
// (18, 21, 'lutff_6/in_3')
// (18, 21, 'lutff_7/in_0')
// (18, 21, 'sp4_h_r_33')
// (18, 21, 'sp4_v_b_29')
// (18, 22, 'local_g1_0')
// (18, 22, 'lutff_2/in_3')
// (18, 22, 'sp4_v_b_16')
// (18, 23, 'local_g0_5')
// (18, 23, 'local_g1_5')
// (18, 23, 'lutff_0/in_3')
// (18, 23, 'lutff_1/in_1')
// (18, 23, 'lutff_2/in_3')
// (18, 23, 'lutff_3/in_0')
// (18, 23, 'lutff_4/in_2')
// (18, 23, 'lutff_5/in_0')
// (18, 23, 'lutff_6/in_3')
// (18, 23, 'lutff_7/in_0')
// (18, 23, 'sp4_h_l_40')
// (18, 23, 'sp4_h_r_21')
// (18, 23, 'sp4_v_b_5')
// (19, 21, 'sp4_h_r_44')
// (19, 23, 'sp4_h_r_32')
// (20, 20, 'sp4_r_v_b_39')
// (20, 21, 'sp4_h_l_44')
// (20, 21, 'sp4_r_v_b_26')
// (20, 22, 'local_g2_7')
// (20, 22, 'lutff_5/in_0')
// (20, 22, 'lutff_6/in_3')
// (20, 22, 'sp4_r_v_b_15')
// (20, 23, 'sp4_h_r_45')
// (20, 23, 'sp4_r_v_b_2')
// (21, 19, 'sp4_v_t_39')
// (21, 20, 'sp4_v_b_39')
// (21, 21, 'sp4_v_b_26')
// (21, 22, 'sp4_v_b_15')
// (21, 23, 'sp4_h_l_45')
// (21, 23, 'sp4_v_b_2')

wire n732;
// (13, 24, 'lutff_7/cout')
// (13, 25, 'carry_in')
// (13, 25, 'carry_in_mux')
// (13, 25, 'lutff_0/in_3')

wire n733;
// (14, 6, 'neigh_op_tnr_0')
// (14, 7, 'neigh_op_rgt_0')
// (14, 8, 'neigh_op_bnr_0')
// (15, 6, 'neigh_op_top_0')
// (15, 7, 'lutff_0/out')
// (15, 8, 'neigh_op_bot_0')
// (16, 6, 'neigh_op_tnl_0')
// (16, 7, 'local_g0_0')
// (16, 7, 'local_g1_0')
// (16, 7, 'lutff_0/in_2')
// (16, 7, 'lutff_0/in_3')
// (16, 7, 'neigh_op_lft_0')
// (16, 8, 'neigh_op_bnl_0')

wire n734;
// (14, 6, 'neigh_op_tnr_1')
// (14, 7, 'local_g1_7')
// (14, 7, 'local_g2_1')
// (14, 7, 'lutff_0/in_0')
// (14, 7, 'lutff_1/in_0')
// (14, 7, 'lutff_2/in_0')
// (14, 7, 'neigh_op_rgt_1')
// (14, 7, 'sp4_h_r_7')
// (14, 8, 'neigh_op_bnr_1')
// (15, 6, 'neigh_op_top_1')
// (15, 7, 'lutff_1/out')
// (15, 7, 'sp4_h_r_18')
// (15, 8, 'neigh_op_bot_1')
// (16, 6, 'neigh_op_tnl_1')
// (16, 7, 'neigh_op_lft_1')
// (16, 7, 'sp4_h_r_31')
// (16, 8, 'neigh_op_bnl_1')
// (17, 7, 'sp4_h_r_42')
// (18, 7, 'sp4_h_l_42')

reg n735 = 0;
// (14, 6, 'neigh_op_tnr_2')
// (14, 7, 'neigh_op_rgt_2')
// (14, 7, 'sp4_r_v_b_36')
// (14, 8, 'neigh_op_bnr_2')
// (14, 8, 'sp4_r_v_b_25')
// (14, 9, 'sp4_r_v_b_12')
// (14, 10, 'sp4_r_v_b_1')
// (15, 6, 'neigh_op_top_2')
// (15, 6, 'sp4_v_t_36')
// (15, 7, 'local_g3_2')
// (15, 7, 'lutff_2/in_3')
// (15, 7, 'lutff_2/out')
// (15, 7, 'sp4_v_b_36')
// (15, 8, 'neigh_op_bot_2')
// (15, 8, 'sp4_v_b_25')
// (15, 9, 'local_g0_4')
// (15, 9, 'lutff_3/in_3')
// (15, 9, 'sp4_v_b_12')
// (15, 10, 'sp4_v_b_1')
// (16, 6, 'neigh_op_tnl_2')
// (16, 7, 'neigh_op_lft_2')
// (16, 8, 'neigh_op_bnl_2')

wire n736;
// (14, 6, 'neigh_op_tnr_3')
// (14, 7, 'neigh_op_rgt_3')
// (14, 8, 'neigh_op_bnr_3')
// (15, 6, 'neigh_op_top_3')
// (15, 7, 'local_g0_3')
// (15, 7, 'lutff_0/in_3')
// (15, 7, 'lutff_3/out')
// (15, 8, 'neigh_op_bot_3')
// (16, 6, 'neigh_op_tnl_3')
// (16, 7, 'neigh_op_lft_3')
// (16, 8, 'neigh_op_bnl_3')

wire n737;
// (14, 6, 'neigh_op_tnr_4')
// (14, 7, 'neigh_op_rgt_4')
// (14, 8, 'neigh_op_bnr_4')
// (15, 6, 'neigh_op_top_4')
// (15, 7, 'local_g0_4')
// (15, 7, 'lutff_4/out')
// (15, 7, 'lutff_7/in_3')
// (15, 8, 'neigh_op_bot_4')
// (16, 6, 'neigh_op_tnl_4')
// (16, 7, 'local_g0_4')
// (16, 7, 'local_g1_4')
// (16, 7, 'lutff_0/in_0')
// (16, 7, 'lutff_1/in_0')
// (16, 7, 'lutff_2/in_0')
// (16, 7, 'neigh_op_lft_4')
// (16, 8, 'neigh_op_bnl_4')

wire n738;
// (14, 6, 'neigh_op_tnr_5')
// (14, 7, 'neigh_op_rgt_5')
// (14, 8, 'neigh_op_bnr_5')
// (15, 6, 'neigh_op_top_5')
// (15, 7, 'local_g3_5')
// (15, 7, 'lutff_1/in_3')
// (15, 7, 'lutff_5/out')
// (15, 8, 'neigh_op_bot_5')
// (16, 6, 'neigh_op_tnl_5')
// (16, 7, 'neigh_op_lft_5')
// (16, 8, 'neigh_op_bnl_5')

wire n739;
// (14, 6, 'neigh_op_tnr_6')
// (14, 7, 'local_g2_6')
// (14, 7, 'local_g3_6')
// (14, 7, 'lutff_0/in_2')
// (14, 7, 'lutff_0/in_3')
// (14, 7, 'neigh_op_rgt_6')
// (14, 8, 'neigh_op_bnr_6')
// (15, 6, 'neigh_op_top_6')
// (15, 7, 'lutff_6/out')
// (15, 8, 'neigh_op_bot_6')
// (16, 6, 'neigh_op_tnl_6')
// (16, 7, 'neigh_op_lft_6')
// (16, 8, 'neigh_op_bnl_6')

reg n740 = 0;
// (14, 6, 'neigh_op_tnr_7')
// (14, 7, 'neigh_op_rgt_7')
// (14, 8, 'neigh_op_bnr_7')
// (15, 2, 'sp12_v_t_22')
// (15, 3, 'sp12_v_b_22')
// (15, 4, 'sp12_v_b_21')
// (15, 5, 'sp12_v_b_18')
// (15, 6, 'neigh_op_top_7')
// (15, 6, 'sp12_v_b_17')
// (15, 7, 'local_g1_7')
// (15, 7, 'lutff_7/in_1')
// (15, 7, 'lutff_7/out')
// (15, 7, 'sp12_v_b_14')
// (15, 8, 'neigh_op_bot_7')
// (15, 8, 'sp12_v_b_13')
// (15, 9, 'sp12_v_b_10')
// (15, 10, 'sp12_v_b_9')
// (15, 11, 'sp12_v_b_6')
// (15, 12, 'local_g3_5')
// (15, 12, 'lutff_5/in_3')
// (15, 12, 'sp12_v_b_5')
// (15, 13, 'sp12_v_b_2')
// (15, 14, 'sp12_v_b_1')
// (16, 6, 'neigh_op_tnl_7')
// (16, 7, 'neigh_op_lft_7')
// (16, 8, 'neigh_op_bnl_7')

wire n741;
// (14, 7, 'lutff_0/cout')
// (14, 7, 'lutff_1/in_3')

wire n742;
// (14, 7, 'lutff_1/cout')
// (14, 7, 'lutff_2/in_3')

wire n743;
// (14, 7, 'lutff_2/cout')
// (14, 7, 'lutff_3/in_3')

wire n744;
// (14, 7, 'lutff_3/cout')
// (14, 7, 'lutff_4/in_3')

wire n745;
// (14, 7, 'lutff_4/cout')
// (14, 7, 'lutff_5/in_3')

reg n746 = 0;
// (14, 8, 'neigh_op_tnr_2')
// (14, 9, 'neigh_op_rgt_2')
// (14, 10, 'neigh_op_bnr_2')
// (15, 8, 'local_g1_2')
// (15, 8, 'lutff_0/in_3')
// (15, 8, 'neigh_op_top_2')
// (15, 9, 'lutff_2/out')
// (15, 10, 'neigh_op_bot_2')
// (16, 8, 'neigh_op_tnl_2')
// (16, 9, 'neigh_op_lft_2')
// (16, 10, 'neigh_op_bnl_2')

reg n747 = 0;
// (14, 8, 'sp4_h_r_1')
// (15, 8, 'local_g1_4')
// (15, 8, 'lutff_7/in_0')
// (15, 8, 'sp4_h_r_12')
// (16, 7, 'neigh_op_tnr_2')
// (16, 8, 'neigh_op_rgt_2')
// (16, 8, 'sp4_h_r_25')
// (16, 9, 'neigh_op_bnr_2')
// (17, 7, 'neigh_op_top_2')
// (17, 8, 'lutff_2/out')
// (17, 8, 'sp4_h_r_36')
// (17, 9, 'neigh_op_bot_2')
// (18, 7, 'neigh_op_tnl_2')
// (18, 8, 'neigh_op_lft_2')
// (18, 8, 'sp4_h_l_36')
// (18, 9, 'neigh_op_bnl_2')

reg n748 = 0;
// (14, 9, 'local_g2_1')
// (14, 9, 'lutff_0/in_1')
// (14, 9, 'neigh_op_tnr_1')
// (14, 10, 'neigh_op_rgt_1')
// (14, 11, 'neigh_op_bnr_1')
// (15, 9, 'neigh_op_top_1')
// (15, 10, 'lutff_1/out')
// (15, 11, 'neigh_op_bot_1')
// (16, 9, 'neigh_op_tnl_1')
// (16, 10, 'neigh_op_lft_1')
// (16, 11, 'neigh_op_bnl_1')

reg n749 = 0;
// (14, 9, 'local_g2_7')
// (14, 9, 'lutff_3/in_0')
// (14, 9, 'neigh_op_tnr_7')
// (14, 10, 'neigh_op_rgt_7')
// (14, 11, 'neigh_op_bnr_7')
// (15, 9, 'neigh_op_top_7')
// (15, 10, 'lutff_7/out')
// (15, 11, 'neigh_op_bot_7')
// (16, 9, 'neigh_op_tnl_7')
// (16, 10, 'neigh_op_lft_7')
// (16, 11, 'neigh_op_bnl_7')

wire n750;
// (14, 9, 'lutff_3/lout')
// (14, 9, 'lutff_4/in_2')

wire n751;
// (14, 9, 'lutff_4/lout')
// (14, 9, 'lutff_5/in_2')

reg n752 = 0;
// (14, 9, 'neigh_op_tnr_0')
// (14, 10, 'neigh_op_rgt_0')
// (14, 11, 'neigh_op_bnr_0')
// (15, 9, 'neigh_op_top_0')
// (15, 10, 'local_g1_0')
// (15, 10, 'lutff_0/out')
// (15, 10, 'lutff_5/in_0')
// (15, 11, 'neigh_op_bot_0')
// (16, 9, 'neigh_op_tnl_0')
// (16, 10, 'neigh_op_lft_0')
// (16, 11, 'neigh_op_bnl_0')

reg n753 = 0;
// (14, 9, 'neigh_op_tnr_4')
// (14, 10, 'neigh_op_rgt_4')
// (14, 10, 'sp4_r_v_b_40')
// (14, 11, 'neigh_op_bnr_4')
// (14, 11, 'sp4_r_v_b_29')
// (14, 12, 'sp4_r_v_b_16')
// (14, 13, 'sp4_r_v_b_5')
// (15, 9, 'neigh_op_top_4')
// (15, 9, 'sp4_v_t_40')
// (15, 10, 'lutff_4/out')
// (15, 10, 'sp4_v_b_40')
// (15, 11, 'neigh_op_bot_4')
// (15, 11, 'sp4_v_b_29')
// (15, 12, 'local_g1_0')
// (15, 12, 'lutff_2/in_3')
// (15, 12, 'sp4_v_b_16')
// (15, 13, 'sp4_v_b_5')
// (16, 9, 'neigh_op_tnl_4')
// (16, 10, 'neigh_op_lft_4')
// (16, 11, 'neigh_op_bnl_4')

reg n754 = 0;
// (14, 9, 'neigh_op_tnr_6')
// (14, 10, 'neigh_op_rgt_6')
// (14, 11, 'neigh_op_bnr_6')
// (15, 9, 'neigh_op_top_6')
// (15, 10, 'local_g2_6')
// (15, 10, 'lutff_0/in_0')
// (15, 10, 'lutff_5/in_1')
// (15, 10, 'lutff_6/out')
// (15, 11, 'neigh_op_bot_6')
// (16, 9, 'neigh_op_tnl_6')
// (16, 10, 'neigh_op_lft_6')
// (16, 11, 'neigh_op_bnl_6')

reg n755 = 0;
// (14, 9, 'sp12_h_r_1')
// (14, 9, 'sp12_v_t_22')
// (14, 10, 'sp12_v_b_22')
// (14, 11, 'sp12_v_b_21')
// (14, 12, 'sp12_v_b_18')
// (14, 13, 'sp12_v_b_17')
// (14, 14, 'sp12_v_b_14')
// (14, 15, 'sp12_v_b_13')
// (14, 16, 'sp12_v_b_10')
// (14, 17, 'sp12_v_b_9')
// (14, 18, 'sp12_v_b_6')
// (14, 19, 'sp12_v_b_5')
// (14, 20, 'sp12_v_b_2')
// (14, 21, 'sp12_h_r_1')
// (14, 21, 'sp12_v_b_1')
// (15, 9, 'sp12_h_r_2')
// (15, 21, 'sp12_h_r_2')
// (16, 9, 'sp12_h_r_5')
// (16, 21, 'sp12_h_r_5')
// (17, 9, 'sp12_h_r_6')
// (17, 21, 'sp12_h_r_6')
// (18, 9, 'local_g1_1')
// (18, 9, 'lutff_1/in_3')
// (18, 9, 'sp12_h_r_9')
// (18, 20, 'neigh_op_tnr_1')
// (18, 21, 'neigh_op_rgt_1')
// (18, 21, 'sp12_h_r_9')
// (18, 22, 'neigh_op_bnr_1')
// (19, 9, 'sp12_h_r_10')
// (19, 20, 'neigh_op_top_1')
// (19, 21, 'lutff_1/out')
// (19, 21, 'sp12_h_r_10')
// (19, 22, 'neigh_op_bot_1')
// (20, 9, 'sp12_h_r_13')
// (20, 20, 'neigh_op_tnl_1')
// (20, 21, 'neigh_op_lft_1')
// (20, 21, 'sp12_h_r_13')
// (20, 22, 'neigh_op_bnl_1')
// (21, 9, 'sp12_h_r_14')
// (21, 21, 'sp12_h_r_14')
// (22, 9, 'sp12_h_r_17')
// (22, 21, 'sp12_h_r_17')
// (23, 9, 'sp12_h_r_18')
// (23, 21, 'sp12_h_r_18')
// (24, 9, 'sp12_h_r_21')
// (24, 21, 'sp12_h_r_21')
// (25, 9, 'sp12_h_r_22')
// (25, 21, 'sp12_h_r_22')
// (26, 9, 'sp12_h_l_22')
// (26, 21, 'sp12_h_l_22')

reg n756 = 0;
// (14, 9, 'sp4_h_r_10')
// (15, 8, 'neigh_op_tnr_1')
// (15, 9, 'neigh_op_rgt_1')
// (15, 9, 'sp4_h_r_23')
// (15, 10, 'neigh_op_bnr_1')
// (16, 8, 'neigh_op_top_1')
// (16, 9, 'lutff_1/out')
// (16, 9, 'sp4_h_r_34')
// (16, 10, 'neigh_op_bot_1')
// (17, 8, 'neigh_op_tnl_1')
// (17, 9, 'neigh_op_lft_1')
// (17, 9, 'sp4_h_r_47')
// (17, 10, 'neigh_op_bnl_1')
// (17, 10, 'sp4_r_v_b_47')
// (17, 11, 'sp4_r_v_b_34')
// (17, 12, 'local_g3_7')
// (17, 12, 'lutff_3/in_3')
// (17, 12, 'sp4_r_v_b_23')
// (17, 13, 'sp4_r_v_b_10')
// (18, 9, 'sp4_h_l_47')
// (18, 9, 'sp4_v_t_47')
// (18, 10, 'sp4_v_b_47')
// (18, 11, 'sp4_v_b_34')
// (18, 12, 'sp4_v_b_23')
// (18, 13, 'sp4_v_b_10')

reg n757 = 0;
// (14, 10, 'local_g0_5')
// (14, 10, 'lutff_4/in_3')
// (14, 10, 'sp4_h_r_5')
// (15, 10, 'sp4_h_r_16')
// (16, 9, 'neigh_op_tnr_4')
// (16, 10, 'neigh_op_rgt_4')
// (16, 10, 'sp4_h_r_29')
// (16, 11, 'neigh_op_bnr_4')
// (17, 9, 'neigh_op_top_4')
// (17, 10, 'lutff_4/out')
// (17, 10, 'sp4_h_r_40')
// (17, 11, 'neigh_op_bot_4')
// (18, 9, 'neigh_op_tnl_4')
// (18, 10, 'neigh_op_lft_4')
// (18, 10, 'sp4_h_l_40')
// (18, 11, 'neigh_op_bnl_4')

reg n758 = 0;
// (14, 10, 'local_g1_1')
// (14, 10, 'lutff_5/in_3')
// (14, 10, 'sp4_h_r_1')
// (15, 10, 'sp4_h_r_12')
// (16, 10, 'sp4_h_r_25')
// (17, 10, 'sp4_h_r_36')
// (17, 11, 'sp4_r_v_b_42')
// (17, 12, 'neigh_op_tnr_1')
// (17, 12, 'sp4_r_v_b_31')
// (17, 13, 'neigh_op_rgt_1')
// (17, 13, 'sp4_r_v_b_18')
// (17, 14, 'neigh_op_bnr_1')
// (17, 14, 'sp4_r_v_b_7')
// (18, 10, 'sp4_h_l_36')
// (18, 10, 'sp4_v_t_42')
// (18, 11, 'sp4_v_b_42')
// (18, 12, 'neigh_op_top_1')
// (18, 12, 'sp4_v_b_31')
// (18, 13, 'lutff_1/out')
// (18, 13, 'sp4_v_b_18')
// (18, 14, 'neigh_op_bot_1')
// (18, 14, 'sp4_v_b_7')
// (19, 12, 'neigh_op_tnl_1')
// (19, 13, 'neigh_op_lft_1')
// (19, 14, 'neigh_op_bnl_1')

reg n759 = 0;
// (14, 10, 'local_g1_3')
// (14, 10, 'lutff_7/in_3')
// (14, 10, 'sp4_h_r_11')
// (15, 10, 'sp4_h_r_22')
// (16, 9, 'neigh_op_tnr_7')
// (16, 10, 'neigh_op_rgt_7')
// (16, 10, 'sp4_h_r_35')
// (16, 11, 'neigh_op_bnr_7')
// (17, 9, 'neigh_op_top_7')
// (17, 10, 'lutff_7/out')
// (17, 10, 'sp4_h_r_46')
// (17, 11, 'neigh_op_bot_7')
// (18, 9, 'neigh_op_tnl_7')
// (18, 10, 'neigh_op_lft_7')
// (18, 10, 'sp4_h_l_46')
// (18, 11, 'neigh_op_bnl_7')

reg n760 = 0;
// (14, 10, 'local_g1_7')
// (14, 10, 'lutff_3/in_3')
// (14, 10, 'sp4_h_r_7')
// (15, 10, 'sp4_h_r_18')
// (16, 9, 'neigh_op_tnr_5')
// (16, 10, 'neigh_op_rgt_5')
// (16, 10, 'sp4_h_r_31')
// (16, 11, 'neigh_op_bnr_5')
// (17, 9, 'neigh_op_top_5')
// (17, 10, 'lutff_5/out')
// (17, 10, 'sp4_h_r_42')
// (17, 11, 'neigh_op_bot_5')
// (18, 9, 'neigh_op_tnl_5')
// (18, 10, 'neigh_op_lft_5')
// (18, 10, 'sp4_h_l_42')
// (18, 11, 'neigh_op_bnl_5')

reg n761 = 0;
// (14, 10, 'neigh_op_tnr_0')
// (14, 10, 'sp4_r_v_b_45')
// (14, 11, 'neigh_op_rgt_0')
// (14, 11, 'sp4_r_v_b_32')
// (14, 12, 'neigh_op_bnr_0')
// (14, 12, 'sp4_r_v_b_21')
// (14, 13, 'sp4_r_v_b_8')
// (15, 9, 'sp4_v_t_45')
// (15, 10, 'neigh_op_top_0')
// (15, 10, 'sp4_v_b_45')
// (15, 11, 'lutff_0/out')
// (15, 11, 'sp4_v_b_32')
// (15, 12, 'local_g0_5')
// (15, 12, 'lutff_4/in_3')
// (15, 12, 'neigh_op_bot_0')
// (15, 12, 'sp4_v_b_21')
// (15, 13, 'sp4_v_b_8')
// (16, 10, 'neigh_op_tnl_0')
// (16, 11, 'neigh_op_lft_0')
// (16, 12, 'neigh_op_bnl_0')

reg n762 = 0;
// (14, 10, 'neigh_op_tnr_1')
// (14, 11, 'neigh_op_rgt_1')
// (14, 12, 'neigh_op_bnr_1')
// (15, 10, 'neigh_op_top_1')
// (15, 11, 'lutff_1/out')
// (15, 12, 'local_g0_1')
// (15, 12, 'lutff_2/in_1')
// (15, 12, 'neigh_op_bot_1')
// (16, 10, 'neigh_op_tnl_1')
// (16, 11, 'neigh_op_lft_1')
// (16, 12, 'neigh_op_bnl_1')

reg n763 = 0;
// (14, 10, 'neigh_op_tnr_4')
// (14, 11, 'neigh_op_rgt_4')
// (14, 12, 'neigh_op_bnr_4')
// (15, 10, 'local_g1_4')
// (15, 10, 'lutff_6/in_3')
// (15, 10, 'neigh_op_top_4')
// (15, 11, 'lutff_4/out')
// (15, 12, 'neigh_op_bot_4')
// (16, 10, 'neigh_op_tnl_4')
// (16, 11, 'neigh_op_lft_4')
// (16, 12, 'neigh_op_bnl_4')

reg n764 = 0;
// (14, 10, 'neigh_op_tnr_5')
// (14, 11, 'neigh_op_rgt_5')
// (14, 12, 'local_g0_5')
// (14, 12, 'lutff_2/in_1')
// (14, 12, 'neigh_op_bnr_5')
// (15, 10, 'neigh_op_top_5')
// (15, 11, 'lutff_5/out')
// (15, 12, 'neigh_op_bot_5')
// (16, 10, 'neigh_op_tnl_5')
// (16, 11, 'neigh_op_lft_5')
// (16, 12, 'neigh_op_bnl_5')

reg n765 = 0;
// (14, 10, 'neigh_op_tnr_6')
// (14, 11, 'neigh_op_rgt_6')
// (14, 12, 'neigh_op_bnr_6')
// (15, 10, 'neigh_op_top_6')
// (15, 11, 'lutff_6/out')
// (15, 12, 'local_g0_6')
// (15, 12, 'lutff_4/in_0')
// (15, 12, 'neigh_op_bot_6')
// (16, 10, 'neigh_op_tnl_6')
// (16, 11, 'neigh_op_lft_6')
// (16, 12, 'neigh_op_bnl_6')

reg n766 = 0;
// (14, 10, 'sp4_r_v_b_43')
// (14, 11, 'sp4_r_v_b_30')
// (14, 12, 'sp4_r_v_b_19')
// (14, 13, 'sp4_r_v_b_6')
// (15, 9, 'sp4_h_r_0')
// (15, 9, 'sp4_v_t_43')
// (15, 10, 'local_g2_3')
// (15, 10, 'lutff_2/in_3')
// (15, 10, 'sp4_v_b_43')
// (15, 11, 'sp4_v_b_30')
// (15, 12, 'sp4_v_b_19')
// (15, 13, 'sp4_v_b_6')
// (16, 8, 'neigh_op_tnr_4')
// (16, 9, 'neigh_op_rgt_4')
// (16, 9, 'sp4_h_r_13')
// (16, 10, 'neigh_op_bnr_4')
// (17, 8, 'neigh_op_top_4')
// (17, 9, 'lutff_4/out')
// (17, 9, 'sp4_h_r_24')
// (17, 10, 'neigh_op_bot_4')
// (18, 8, 'neigh_op_tnl_4')
// (18, 9, 'neigh_op_lft_4')
// (18, 9, 'sp4_h_r_37')
// (18, 10, 'neigh_op_bnl_4')
// (19, 9, 'sp4_h_l_37')

wire n767;
// (14, 11, 'neigh_op_tnr_2')
// (14, 12, 'local_g2_2')
// (14, 12, 'lutff_3/in_3')
// (14, 12, 'neigh_op_rgt_2')
// (14, 13, 'neigh_op_bnr_2')
// (15, 11, 'neigh_op_top_2')
// (15, 12, 'lutff_2/out')
// (15, 13, 'neigh_op_bot_2')
// (16, 11, 'neigh_op_tnl_2')
// (16, 12, 'neigh_op_lft_2')
// (16, 13, 'neigh_op_bnl_2')

wire n768;
// (14, 11, 'neigh_op_tnr_4')
// (14, 12, 'local_g2_4')
// (14, 12, 'lutff_3/in_1')
// (14, 12, 'neigh_op_rgt_4')
// (14, 13, 'neigh_op_bnr_4')
// (15, 11, 'neigh_op_top_4')
// (15, 12, 'lutff_4/out')
// (15, 13, 'neigh_op_bot_4')
// (16, 11, 'neigh_op_tnl_4')
// (16, 12, 'neigh_op_lft_4')
// (16, 13, 'neigh_op_bnl_4')

wire n769;
// (14, 11, 'sp4_r_v_b_37')
// (14, 12, 'local_g0_0')
// (14, 12, 'lutff_5/in_1')
// (14, 12, 'sp4_r_v_b_24')
// (14, 13, 'neigh_op_tnr_0')
// (14, 13, 'sp4_r_v_b_13')
// (14, 14, 'neigh_op_rgt_0')
// (14, 14, 'sp4_r_v_b_0')
// (14, 15, 'neigh_op_bnr_0')
// (15, 10, 'sp4_v_t_37')
// (15, 11, 'sp4_v_b_37')
// (15, 12, 'local_g3_0')
// (15, 12, 'lutff_0/in_3')
// (15, 12, 'sp4_v_b_24')
// (15, 13, 'neigh_op_top_0')
// (15, 13, 'sp4_r_v_b_44')
// (15, 13, 'sp4_v_b_13')
// (15, 14, 'lutff_0/out')
// (15, 14, 'sp4_r_v_b_33')
// (15, 14, 'sp4_v_b_0')
// (15, 15, 'neigh_op_bot_0')
// (15, 15, 'sp4_r_v_b_20')
// (15, 16, 'sp4_r_v_b_9')
// (16, 12, 'sp4_h_r_9')
// (16, 12, 'sp4_v_t_44')
// (16, 13, 'neigh_op_tnl_0')
// (16, 13, 'sp4_v_b_44')
// (16, 14, 'neigh_op_lft_0')
// (16, 14, 'sp4_v_b_33')
// (16, 15, 'local_g2_0')
// (16, 15, 'lutff_7/in_3')
// (16, 15, 'neigh_op_bnl_0')
// (16, 15, 'sp4_v_b_20')
// (16, 16, 'sp4_v_b_9')
// (17, 12, 'sp4_h_r_20')
// (18, 12, 'sp4_h_r_33')
// (19, 12, 'local_g3_4')
// (19, 12, 'lutff_4/in_3')
// (19, 12, 'sp4_h_r_44')
// (20, 12, 'sp4_h_l_44')

reg n770 = 0;
// (14, 11, 'sp4_r_v_b_45')
// (14, 12, 'local_g0_3')
// (14, 12, 'lutff_4/in_3')
// (14, 12, 'lutff_6/in_3')
// (14, 12, 'sp4_r_v_b_32')
// (14, 13, 'neigh_op_tnr_4')
// (14, 13, 'sp4_r_v_b_21')
// (14, 14, 'local_g3_4')
// (14, 14, 'lutff_0/in_3')
// (14, 14, 'neigh_op_rgt_4')
// (14, 14, 'sp4_r_v_b_8')
// (14, 15, 'local_g1_4')
// (14, 15, 'lutff_7/in_0')
// (14, 15, 'neigh_op_bnr_4')
// (15, 10, 'sp4_v_t_45')
// (15, 11, 'sp4_r_v_b_44')
// (15, 11, 'sp4_v_b_45')
// (15, 12, 'sp4_r_v_b_33')
// (15, 12, 'sp4_v_b_32')
// (15, 13, 'local_g1_4')
// (15, 13, 'lutff_6/in_3')
// (15, 13, 'lutff_7/in_0')
// (15, 13, 'neigh_op_top_4')
// (15, 13, 'sp4_r_v_b_20')
// (15, 13, 'sp4_v_b_21')
// (15, 14, 'local_g1_4')
// (15, 14, 'lutff_3/in_2')
// (15, 14, 'lutff_4/in_1')
// (15, 14, 'lutff_4/out')
// (15, 14, 'lutff_5/in_2')
// (15, 14, 'lutff_6/in_1')
// (15, 14, 'sp4_r_v_b_9')
// (15, 14, 'sp4_v_b_8')
// (15, 15, 'neigh_op_bot_4')
// (16, 10, 'sp4_v_t_44')
// (16, 11, 'sp4_v_b_44')
// (16, 12, 'local_g3_1')
// (16, 12, 'lutff_1/in_3')
// (16, 12, 'lutff_5/in_3')
// (16, 12, 'sp4_v_b_33')
// (16, 13, 'local_g2_4')
// (16, 13, 'lutff_1/in_3')
// (16, 13, 'lutff_3/in_3')
// (16, 13, 'neigh_op_tnl_4')
// (16, 13, 'sp4_v_b_20')
// (16, 14, 'local_g0_4')
// (16, 14, 'lutff_3/in_3')
// (16, 14, 'neigh_op_lft_4')
// (16, 14, 'sp4_v_b_9')
// (16, 15, 'neigh_op_bnl_4')

reg n771 = 0;
// (14, 11, 'sp4_r_v_b_47')
// (14, 12, 'local_g0_1')
// (14, 12, 'lutff_4/in_1')
// (14, 12, 'sp4_r_v_b_34')
// (14, 13, 'neigh_op_tnr_5')
// (14, 13, 'sp4_r_v_b_23')
// (14, 14, 'neigh_op_rgt_5')
// (14, 14, 'sp4_r_v_b_10')
// (14, 15, 'local_g1_5')
// (14, 15, 'lutff_6/in_0')
// (14, 15, 'lutff_7/in_1')
// (14, 15, 'neigh_op_bnr_5')
// (15, 10, 'sp4_v_t_47')
// (15, 11, 'sp4_v_b_47')
// (15, 12, 'sp4_v_b_34')
// (15, 13, 'neigh_op_top_5')
// (15, 13, 'sp4_v_b_23')
// (15, 14, 'local_g2_5')
// (15, 14, 'lutff_3/in_0')
// (15, 14, 'lutff_4/in_3')
// (15, 14, 'lutff_5/in_0')
// (15, 14, 'lutff_5/out')
// (15, 14, 'lutff_6/in_3')
// (15, 14, 'sp4_v_b_10')
// (15, 15, 'neigh_op_bot_5')
// (16, 13, 'neigh_op_tnl_5')
// (16, 14, 'neigh_op_lft_5')
// (16, 15, 'neigh_op_bnl_5')

wire n772;
// (14, 12, 'lutff_0/lout')
// (14, 12, 'lutff_1/in_2')

wire n773;
// (14, 12, 'lutff_4/lout')
// (14, 12, 'lutff_5/in_2')

wire n774;
// (14, 12, 'lutff_5/lout')
// (14, 12, 'lutff_6/in_2')

wire n775;
// (14, 12, 'neigh_op_tnr_1')
// (14, 13, 'neigh_op_rgt_1')
// (14, 14, 'neigh_op_bnr_1')
// (15, 12, 'neigh_op_top_1')
// (15, 13, 'local_g2_1')
// (15, 13, 'lutff_1/out')
// (15, 13, 'lutff_3/in_2')
// (15, 14, 'neigh_op_bot_1')
// (16, 12, 'neigh_op_tnl_1')
// (16, 13, 'neigh_op_lft_1')
// (16, 14, 'neigh_op_bnl_1')

wire n776;
// (14, 12, 'neigh_op_tnr_4')
// (14, 13, 'neigh_op_rgt_4')
// (14, 14, 'neigh_op_bnr_4')
// (15, 12, 'neigh_op_top_4')
// (15, 13, 'lutff_4/out')
// (15, 14, 'local_g0_4')
// (15, 14, 'lutff_0/in_2')
// (15, 14, 'lutff_3/in_1')
// (15, 14, 'neigh_op_bot_4')
// (16, 12, 'local_g2_4')
// (16, 12, 'lutff_7/in_3')
// (16, 12, 'neigh_op_tnl_4')
// (16, 13, 'neigh_op_lft_4')
// (16, 14, 'neigh_op_bnl_4')

wire n777;
// (14, 12, 'neigh_op_tnr_5')
// (14, 13, 'neigh_op_rgt_5')
// (14, 13, 'sp4_r_v_b_42')
// (14, 14, 'neigh_op_bnr_5')
// (14, 14, 'sp4_r_v_b_31')
// (14, 15, 'sp4_r_v_b_18')
// (14, 16, 'sp4_r_v_b_7')
// (15, 12, 'neigh_op_top_5')
// (15, 12, 'sp4_v_t_42')
// (15, 13, 'local_g2_5')
// (15, 13, 'lutff_2/in_1')
// (15, 13, 'lutff_3/in_0')
// (15, 13, 'lutff_5/out')
// (15, 13, 'sp4_v_b_42')
// (15, 14, 'neigh_op_bot_5')
// (15, 14, 'sp4_v_b_31')
// (15, 15, 'sp4_v_b_18')
// (15, 16, 'local_g1_7')
// (15, 16, 'lutff_3/in_1')
// (15, 16, 'sp4_v_b_7')
// (16, 12, 'neigh_op_tnl_5')
// (16, 13, 'neigh_op_lft_5')
// (16, 14, 'neigh_op_bnl_5')

reg n778 = 0;
// (14, 12, 'neigh_op_tnr_6')
// (14, 12, 'sp4_r_v_b_41')
// (14, 13, 'neigh_op_rgt_6')
// (14, 13, 'sp4_r_v_b_28')
// (14, 14, 'neigh_op_bnr_6')
// (14, 14, 'sp4_r_v_b_17')
// (14, 15, 'sp4_r_v_b_4')
// (15, 11, 'sp4_v_t_41')
// (15, 12, 'neigh_op_top_6')
// (15, 12, 'sp4_v_b_41')
// (15, 13, 'local_g3_6')
// (15, 13, 'lutff_0/in_3')
// (15, 13, 'lutff_4/in_3')
// (15, 13, 'lutff_6/out')
// (15, 13, 'sp4_r_v_b_45')
// (15, 13, 'sp4_v_b_28')
// (15, 14, 'neigh_op_bot_6')
// (15, 14, 'sp4_r_v_b_32')
// (15, 14, 'sp4_v_b_17')
// (15, 15, 'sp4_h_r_10')
// (15, 15, 'sp4_r_v_b_21')
// (15, 15, 'sp4_v_b_4')
// (15, 16, 'sp4_r_v_b_8')
// (16, 12, 'local_g3_6')
// (16, 12, 'lutff_2/in_3')
// (16, 12, 'neigh_op_tnl_6')
// (16, 12, 'sp4_v_t_45')
// (16, 13, 'neigh_op_lft_6')
// (16, 13, 'sp4_v_b_45')
// (16, 14, 'local_g2_6')
// (16, 14, 'local_g3_6')
// (16, 14, 'lutff_0/in_3')
// (16, 14, 'lutff_1/in_2')
// (16, 14, 'lutff_5/in_1')
// (16, 14, 'neigh_op_bnl_6')
// (16, 14, 'sp4_v_b_32')
// (16, 15, 'local_g0_5')
// (16, 15, 'lutff_0/in_3')
// (16, 15, 'lutff_3/in_0')
// (16, 15, 'sp4_h_r_23')
// (16, 15, 'sp4_v_b_21')
// (16, 16, 'sp4_v_b_8')
// (17, 15, 'sp4_h_r_34')
// (18, 15, 'local_g2_7')
// (18, 15, 'lutff_0/in_1')
// (18, 15, 'sp4_h_r_47')
// (19, 15, 'sp4_h_l_47')

reg n779 = 0;
// (14, 12, 'neigh_op_tnr_7')
// (14, 13, 'neigh_op_rgt_7')
// (14, 14, 'neigh_op_bnr_7')
// (15, 12, 'neigh_op_top_7')
// (15, 13, 'local_g1_7')
// (15, 13, 'lutff_1/in_3')
// (15, 13, 'lutff_4/in_0')
// (15, 13, 'lutff_7/out')
// (15, 14, 'local_g1_7')
// (15, 14, 'lutff_7/in_1')
// (15, 14, 'neigh_op_bot_7')
// (16, 12, 'local_g3_7')
// (16, 12, 'lutff_2/in_0')
// (16, 12, 'neigh_op_tnl_7')
// (16, 13, 'neigh_op_lft_7')
// (16, 14, 'neigh_op_bnl_7')

wire n780;
// (14, 12, 'sp4_r_v_b_38')
// (14, 13, 'neigh_op_tnr_7')
// (14, 13, 'sp4_r_v_b_27')
// (14, 14, 'neigh_op_rgt_7')
// (14, 14, 'sp4_r_v_b_14')
// (14, 15, 'neigh_op_bnr_7')
// (14, 15, 'sp4_r_v_b_3')
// (15, 11, 'sp4_v_t_38')
// (15, 12, 'sp4_v_b_38')
// (15, 13, 'neigh_op_top_7')
// (15, 13, 'sp4_v_b_27')
// (15, 14, 'lutff_7/out')
// (15, 14, 'sp4_v_b_14')
// (15, 15, 'neigh_op_bot_7')
// (15, 15, 'sp4_h_r_3')
// (15, 15, 'sp4_v_b_3')
// (16, 13, 'neigh_op_tnl_7')
// (16, 14, 'local_g1_7')
// (16, 14, 'lutff_0/in_0')
// (16, 14, 'lutff_1/in_3')
// (16, 14, 'lutff_5/in_3')
// (16, 14, 'neigh_op_lft_7')
// (16, 15, 'local_g3_7')
// (16, 15, 'lutff_0/in_0')
// (16, 15, 'lutff_3/in_3')
// (16, 15, 'neigh_op_bnl_7')
// (16, 15, 'sp4_h_r_14')
// (17, 15, 'sp4_h_r_27')
// (18, 15, 'local_g3_6')
// (18, 15, 'lutff_0/in_3')
// (18, 15, 'sp4_h_r_38')
// (19, 15, 'sp4_h_l_38')

wire n781;
// (14, 13, 'neigh_op_tnr_1')
// (14, 14, 'neigh_op_rgt_1')
// (14, 15, 'neigh_op_bnr_1')
// (15, 13, 'neigh_op_top_1')
// (15, 13, 'sp4_r_v_b_46')
// (15, 14, 'lutff_1/out')
// (15, 14, 'sp4_r_v_b_35')
// (15, 15, 'neigh_op_bot_1')
// (15, 15, 'sp4_r_v_b_22')
// (15, 16, 'local_g2_3')
// (15, 16, 'lutff_3/in_0')
// (15, 16, 'sp4_r_v_b_11')
// (15, 17, 'sp4_r_v_b_39')
// (15, 18, 'sp4_r_v_b_26')
// (15, 19, 'sp4_r_v_b_15')
// (15, 20, 'sp4_r_v_b_2')
// (16, 12, 'sp4_v_t_46')
// (16, 13, 'neigh_op_tnl_1')
// (16, 13, 'sp4_v_b_46')
// (16, 14, 'neigh_op_lft_1')
// (16, 14, 'sp4_v_b_35')
// (16, 15, 'neigh_op_bnl_1')
// (16, 15, 'sp4_v_b_22')
// (16, 16, 'sp4_v_b_11')
// (16, 16, 'sp4_v_t_39')
// (16, 17, 'sp4_v_b_39')
// (16, 18, 'sp4_v_b_26')
// (16, 19, 'sp4_v_b_15')
// (16, 20, 'local_g1_2')
// (16, 20, 'lutff_6/in_3')
// (16, 20, 'sp4_v_b_2')

wire n782;
// (14, 13, 'neigh_op_tnr_6')
// (14, 14, 'neigh_op_rgt_6')
// (14, 14, 'sp4_h_r_1')
// (14, 15, 'neigh_op_bnr_6')
// (15, 12, 'sp4_r_v_b_37')
// (15, 13, 'local_g0_6')
// (15, 13, 'local_g1_6')
// (15, 13, 'lutff_2/in_3')
// (15, 13, 'lutff_3/in_1')
// (15, 13, 'neigh_op_top_6')
// (15, 13, 'sp4_r_v_b_24')
// (15, 14, 'local_g3_6')
// (15, 14, 'lutff_0/in_3')
// (15, 14, 'lutff_6/out')
// (15, 14, 'sp4_h_r_12')
// (15, 14, 'sp4_r_v_b_13')
// (15, 15, 'neigh_op_bot_6')
// (15, 15, 'sp4_r_v_b_0')
// (16, 11, 'sp4_v_t_37')
// (16, 12, 'local_g3_5')
// (16, 12, 'lutff_4/in_0')
// (16, 12, 'sp4_v_b_37')
// (16, 13, 'neigh_op_tnl_6')
// (16, 13, 'sp4_v_b_24')
// (16, 14, 'neigh_op_lft_6')
// (16, 14, 'sp4_h_r_25')
// (16, 14, 'sp4_v_b_13')
// (16, 15, 'neigh_op_bnl_6')
// (16, 15, 'sp4_v_b_0')
// (17, 14, 'sp4_h_r_36')
// (17, 15, 'sp4_r_v_b_43')
// (17, 16, 'sp4_r_v_b_30')
// (17, 17, 'sp4_r_v_b_19')
// (17, 18, 'sp4_r_v_b_6')
// (18, 14, 'sp4_h_l_36')
// (18, 14, 'sp4_v_t_43')
// (18, 15, 'sp4_v_b_43')
// (18, 16, 'sp4_v_b_30')
// (18, 17, 'sp4_v_b_19')
// (18, 18, 'sp4_h_r_6')
// (18, 18, 'sp4_v_b_6')
// (19, 18, 'sp4_h_r_19')
// (20, 18, 'local_g3_6')
// (20, 18, 'lutff_2/in_3')
// (20, 18, 'sp4_h_r_30')
// (21, 18, 'sp4_h_r_43')
// (22, 18, 'sp4_h_l_43')

reg n783 = 0;
// (14, 13, 'sp4_h_r_11')
// (15, 13, 'sp4_h_r_22')
// (16, 13, 'sp4_h_r_35')
// (17, 13, 'local_g2_6')
// (17, 13, 'lutff_1/in_3')
// (17, 13, 'sp4_h_r_46')
// (18, 13, 'sp4_h_l_46')
// (18, 13, 'sp4_h_r_3')
// (19, 13, 'sp4_h_r_14')
// (20, 13, 'sp4_h_r_27')
// (21, 13, 'neigh_op_tnr_6')
// (21, 13, 'sp4_h_r_38')
// (21, 14, 'neigh_op_rgt_6')
// (21, 14, 'sp4_r_v_b_44')
// (21, 15, 'neigh_op_bnr_6')
// (21, 15, 'sp4_r_v_b_33')
// (21, 16, 'sp4_r_v_b_20')
// (21, 17, 'sp4_r_v_b_9')
// (22, 13, 'neigh_op_top_6')
// (22, 13, 'sp4_h_l_38')
// (22, 13, 'sp4_v_t_44')
// (22, 14, 'lutff_6/out')
// (22, 14, 'sp4_v_b_44')
// (22, 15, 'neigh_op_bot_6')
// (22, 15, 'sp4_v_b_33')
// (22, 16, 'sp4_v_b_20')
// (22, 17, 'sp4_v_b_9')
// (23, 13, 'neigh_op_tnl_6')
// (23, 14, 'neigh_op_lft_6')
// (23, 15, 'neigh_op_bnl_6')

reg n784 = 0;
// (14, 13, 'sp4_h_r_2')
// (15, 13, 'sp4_h_r_15')
// (16, 13, 'sp4_h_r_26')
// (17, 13, 'local_g3_7')
// (17, 13, 'lutff_5/in_3')
// (17, 13, 'sp4_h_r_39')
// (18, 13, 'sp4_h_l_39')
// (18, 13, 'sp4_h_r_11')
// (19, 13, 'sp4_h_r_22')
// (20, 13, 'sp4_h_r_35')
// (21, 13, 'neigh_op_tnr_7')
// (21, 13, 'sp4_h_r_46')
// (21, 14, 'neigh_op_rgt_7')
// (21, 14, 'sp4_r_v_b_46')
// (21, 15, 'neigh_op_bnr_7')
// (21, 15, 'sp4_r_v_b_35')
// (21, 16, 'sp4_r_v_b_22')
// (21, 17, 'sp4_r_v_b_11')
// (22, 13, 'neigh_op_top_7')
// (22, 13, 'sp4_h_l_46')
// (22, 13, 'sp4_v_t_46')
// (22, 14, 'lutff_7/out')
// (22, 14, 'sp4_v_b_46')
// (22, 15, 'neigh_op_bot_7')
// (22, 15, 'sp4_v_b_35')
// (22, 16, 'sp4_v_b_22')
// (22, 17, 'sp4_v_b_11')
// (23, 13, 'neigh_op_tnl_7')
// (23, 14, 'neigh_op_lft_7')
// (23, 15, 'neigh_op_bnl_7')

reg n785 = 0;
// (14, 13, 'sp4_r_v_b_46')
// (14, 14, 'neigh_op_tnr_3')
// (14, 14, 'sp4_r_v_b_35')
// (14, 15, 'neigh_op_rgt_3')
// (14, 15, 'sp4_r_v_b_22')
// (14, 16, 'neigh_op_bnr_3')
// (14, 16, 'sp4_r_v_b_11')
// (15, 12, 'sp4_v_t_46')
// (15, 13, 'sp4_v_b_46')
// (15, 14, 'neigh_op_top_3')
// (15, 14, 'sp4_v_b_35')
// (15, 15, 'lutff_3/out')
// (15, 15, 'sp4_v_b_22')
// (15, 16, 'neigh_op_bot_3')
// (15, 16, 'sp4_h_r_5')
// (15, 16, 'sp4_v_b_11')
// (16, 14, 'neigh_op_tnl_3')
// (16, 15, 'neigh_op_lft_3')
// (16, 16, 'neigh_op_bnl_3')
// (16, 16, 'sp4_h_r_16')
// (17, 16, 'sp4_h_r_29')
// (18, 16, 'sp4_h_r_40')
// (19, 16, 'sp4_h_l_40')
// (19, 16, 'sp4_h_r_5')
// (20, 16, 'sp4_h_r_16')
// (21, 16, 'local_g2_5')
// (21, 16, 'lutff_4/in_1')
// (21, 16, 'sp4_h_r_29')
// (22, 16, 'sp4_h_r_40')
// (23, 16, 'sp4_h_l_40')

reg n786 = 0;
// (14, 14, 'neigh_op_tnr_1')
// (14, 15, 'neigh_op_rgt_1')
// (14, 16, 'neigh_op_bnr_1')
// (15, 14, 'neigh_op_top_1')
// (15, 14, 'sp4_r_v_b_46')
// (15, 15, 'lutff_1/out')
// (15, 15, 'sp4_r_v_b_35')
// (15, 16, 'neigh_op_bot_1')
// (15, 16, 'sp4_r_v_b_22')
// (15, 17, 'sp4_r_v_b_11')
// (16, 13, 'sp4_h_r_4')
// (16, 13, 'sp4_v_t_46')
// (16, 14, 'neigh_op_tnl_1')
// (16, 14, 'sp4_v_b_46')
// (16, 15, 'neigh_op_lft_1')
// (16, 15, 'sp4_v_b_35')
// (16, 16, 'neigh_op_bnl_1')
// (16, 16, 'sp4_v_b_22')
// (16, 17, 'sp4_v_b_11')
// (17, 13, 'sp4_h_r_17')
// (18, 13, 'sp4_h_r_28')
// (19, 13, 'local_g2_1')
// (19, 13, 'lutff_2/in_1')
// (19, 13, 'sp4_h_r_41')
// (20, 13, 'sp4_h_l_41')

reg n787 = 0;
// (14, 14, 'neigh_op_tnr_2')
// (14, 15, 'neigh_op_rgt_2')
// (14, 15, 'sp4_h_r_9')
// (14, 16, 'neigh_op_bnr_2')
// (15, 14, 'neigh_op_top_2')
// (15, 15, 'lutff_2/out')
// (15, 15, 'sp4_h_r_20')
// (15, 16, 'neigh_op_bot_2')
// (16, 14, 'neigh_op_tnl_2')
// (16, 15, 'neigh_op_lft_2')
// (16, 15, 'sp4_h_r_33')
// (16, 16, 'neigh_op_bnl_2')
// (17, 15, 'sp4_h_r_44')
// (18, 15, 'sp4_h_l_44')
// (18, 15, 'sp4_h_r_0')
// (19, 15, 'sp4_h_r_13')
// (20, 15, 'sp4_h_r_24')
// (21, 12, 'sp4_r_v_b_37')
// (21, 13, 'local_g1_0')
// (21, 13, 'lutff_6/in_1')
// (21, 13, 'sp4_r_v_b_24')
// (21, 14, 'sp4_r_v_b_13')
// (21, 15, 'sp4_h_r_37')
// (21, 15, 'sp4_r_v_b_0')
// (22, 11, 'sp4_v_t_37')
// (22, 12, 'sp4_v_b_37')
// (22, 13, 'sp4_v_b_24')
// (22, 14, 'sp4_v_b_13')
// (22, 15, 'sp4_h_l_37')
// (22, 15, 'sp4_v_b_0')

reg n788 = 0;
// (14, 14, 'neigh_op_tnr_4')
// (14, 15, 'neigh_op_rgt_4')
// (14, 16, 'neigh_op_bnr_4')
// (15, 14, 'neigh_op_top_4')
// (15, 15, 'lutff_4/out')
// (15, 15, 'sp4_h_r_8')
// (15, 16, 'neigh_op_bot_4')
// (16, 14, 'neigh_op_tnl_4')
// (16, 15, 'neigh_op_lft_4')
// (16, 15, 'sp4_h_r_21')
// (16, 16, 'neigh_op_bnl_4')
// (17, 15, 'sp4_h_r_32')
// (18, 15, 'sp4_h_r_45')
// (19, 15, 'sp4_h_l_45')
// (19, 15, 'sp4_h_r_4')
// (20, 15, 'sp4_h_r_17')
// (21, 15, 'sp4_h_r_28')
// (22, 15, 'sp4_h_r_41')
// (22, 16, 'local_g3_4')
// (22, 16, 'lutff_6/in_1')
// (22, 16, 'sp4_r_v_b_44')
// (22, 17, 'sp4_r_v_b_33')
// (22, 18, 'sp4_r_v_b_20')
// (22, 19, 'sp4_r_v_b_9')
// (23, 15, 'sp4_h_l_41')
// (23, 15, 'sp4_v_t_44')
// (23, 16, 'sp4_v_b_44')
// (23, 17, 'sp4_v_b_33')
// (23, 18, 'sp4_v_b_20')
// (23, 19, 'sp4_v_b_9')

reg n789 = 0;
// (14, 14, 'neigh_op_tnr_5')
// (14, 15, 'neigh_op_rgt_5')
// (14, 16, 'neigh_op_bnr_5')
// (15, 14, 'neigh_op_top_5')
// (15, 15, 'lutff_5/out')
// (15, 15, 'sp4_r_v_b_43')
// (15, 16, 'neigh_op_bot_5')
// (15, 16, 'sp4_r_v_b_30')
// (15, 17, 'sp4_r_v_b_19')
// (15, 18, 'sp4_r_v_b_6')
// (16, 14, 'neigh_op_tnl_5')
// (16, 14, 'sp4_v_t_43')
// (16, 15, 'neigh_op_lft_5')
// (16, 15, 'sp4_v_b_43')
// (16, 16, 'neigh_op_bnl_5')
// (16, 16, 'sp4_v_b_30')
// (16, 17, 'sp4_v_b_19')
// (16, 18, 'sp4_h_r_0')
// (16, 18, 'sp4_v_b_6')
// (17, 18, 'sp4_h_r_13')
// (18, 18, 'sp4_h_r_24')
// (19, 18, 'local_g2_5')
// (19, 18, 'lutff_4/in_1')
// (19, 18, 'sp4_h_r_37')
// (20, 18, 'sp4_h_l_37')

reg n790 = 0;
// (14, 14, 'neigh_op_tnr_6')
// (14, 15, 'neigh_op_rgt_6')
// (14, 15, 'sp4_r_v_b_44')
// (14, 16, 'neigh_op_bnr_6')
// (14, 16, 'sp4_r_v_b_33')
// (14, 17, 'sp4_r_v_b_20')
// (14, 18, 'sp4_r_v_b_9')
// (15, 14, 'neigh_op_top_6')
// (15, 14, 'sp4_h_r_2')
// (15, 14, 'sp4_v_t_44')
// (15, 15, 'lutff_6/out')
// (15, 15, 'sp4_v_b_44')
// (15, 16, 'neigh_op_bot_6')
// (15, 16, 'sp4_v_b_33')
// (15, 17, 'sp4_v_b_20')
// (15, 18, 'sp4_v_b_9')
// (16, 14, 'neigh_op_tnl_6')
// (16, 14, 'sp4_h_r_15')
// (16, 15, 'neigh_op_lft_6')
// (16, 16, 'neigh_op_bnl_6')
// (17, 14, 'sp4_h_r_26')
// (18, 14, 'sp4_h_r_39')
// (19, 14, 'local_g1_2')
// (19, 14, 'lutff_4/in_1')
// (19, 14, 'sp4_h_l_39')
// (19, 14, 'sp4_h_r_2')
// (20, 14, 'sp4_h_r_15')
// (21, 14, 'sp4_h_r_26')
// (22, 14, 'sp4_h_r_39')
// (23, 14, 'sp4_h_l_39')

reg n791 = 0;
// (14, 14, 'neigh_op_tnr_7')
// (14, 15, 'neigh_op_rgt_7')
// (14, 15, 'sp4_r_v_b_46')
// (14, 16, 'neigh_op_bnr_7')
// (14, 16, 'sp4_r_v_b_35')
// (14, 17, 'sp4_r_v_b_22')
// (14, 18, 'sp4_r_v_b_11')
// (15, 14, 'neigh_op_top_7')
// (15, 14, 'sp4_h_r_11')
// (15, 14, 'sp4_v_t_46')
// (15, 15, 'lutff_7/out')
// (15, 15, 'sp4_v_b_46')
// (15, 16, 'neigh_op_bot_7')
// (15, 16, 'sp4_v_b_35')
// (15, 17, 'sp4_v_b_22')
// (15, 18, 'sp4_v_b_11')
// (16, 14, 'neigh_op_tnl_7')
// (16, 14, 'sp4_h_r_22')
// (16, 15, 'neigh_op_lft_7')
// (16, 16, 'neigh_op_bnl_7')
// (17, 14, 'local_g3_3')
// (17, 14, 'lutff_7/in_1')
// (17, 14, 'sp4_h_r_35')
// (18, 14, 'sp4_h_r_46')
// (19, 14, 'sp4_h_l_46')

reg n792 = 0;
// (14, 14, 'sp12_h_r_0')
// (15, 14, 'sp12_h_r_3')
// (16, 14, 'sp12_h_r_4')
// (17, 14, 'sp12_h_r_7')
// (18, 14, 'sp12_h_r_8')
// (19, 14, 'local_g1_3')
// (19, 14, 'lutff_3/in_3')
// (19, 14, 'sp12_h_r_11')
// (20, 14, 'sp12_h_r_12')
// (21, 14, 'sp12_h_r_15')
// (22, 14, 'sp12_h_r_16')
// (23, 13, 'neigh_op_tnr_6')
// (23, 14, 'neigh_op_rgt_6')
// (23, 14, 'sp12_h_r_19')
// (23, 15, 'neigh_op_bnr_6')
// (24, 13, 'neigh_op_top_6')
// (24, 14, 'lutff_6/out')
// (24, 14, 'sp12_h_r_20')
// (24, 15, 'neigh_op_bot_6')
// (25, 13, 'neigh_op_tnl_6')
// (25, 14, 'neigh_op_lft_6')
// (25, 14, 'sp12_h_r_23')
// (25, 15, 'neigh_op_bnl_6')
// (26, 14, 'sp12_h_l_23')

wire n793;
// (14, 14, 'sp4_r_v_b_42')
// (14, 15, 'neigh_op_tnr_1')
// (14, 15, 'sp4_r_v_b_31')
// (14, 16, 'neigh_op_rgt_1')
// (14, 16, 'sp4_r_v_b_18')
// (14, 17, 'neigh_op_bnr_1')
// (14, 17, 'sp4_r_v_b_7')
// (15, 13, 'sp4_v_t_42')
// (15, 14, 'sp4_v_b_42')
// (15, 15, 'neigh_op_top_1')
// (15, 15, 'sp4_v_b_31')
// (15, 16, 'lutff_1/out')
// (15, 16, 'sp4_v_b_18')
// (15, 17, 'neigh_op_bot_1')
// (15, 17, 'sp4_h_r_7')
// (15, 17, 'sp4_v_b_7')
// (16, 15, 'neigh_op_tnl_1')
// (16, 16, 'neigh_op_lft_1')
// (16, 17, 'neigh_op_bnl_1')
// (16, 17, 'sp4_h_r_18')
// (17, 17, 'sp4_h_r_31')
// (18, 17, 'sp4_h_r_42')
// (19, 17, 'sp4_h_l_42')
// (19, 17, 'sp4_h_r_10')
// (19, 17, 'sp4_h_r_7')
// (20, 17, 'local_g0_2')
// (20, 17, 'lutff_global/cen')
// (20, 17, 'sp4_h_r_18')
// (20, 17, 'sp4_h_r_23')
// (21, 17, 'sp4_h_r_31')
// (21, 17, 'sp4_h_r_34')
// (22, 14, 'sp4_r_v_b_47')
// (22, 15, 'sp4_r_v_b_34')
// (22, 16, 'sp4_r_v_b_23')
// (22, 17, 'sp4_h_r_42')
// (22, 17, 'sp4_h_r_47')
// (22, 17, 'sp4_r_v_b_10')
// (22, 18, 'sp4_r_v_b_47')
// (22, 19, 'sp4_r_v_b_34')
// (22, 20, 'sp4_r_v_b_23')
// (22, 21, 'sp4_r_v_b_10')
// (22, 22, 'sp4_r_v_b_43')
// (22, 23, 'sp4_r_v_b_30')
// (22, 24, 'sp4_r_v_b_19')
// (22, 25, 'sp4_r_v_b_6')
// (23, 13, 'local_g0_2')
// (23, 13, 'lutff_global/cen')
// (23, 13, 'sp4_h_r_10')
// (23, 13, 'sp4_v_t_47')
// (23, 14, 'sp4_v_b_47')
// (23, 15, 'sp4_v_b_34')
// (23, 16, 'sp4_v_b_23')
// (23, 17, 'sp4_h_l_42')
// (23, 17, 'sp4_h_l_47')
// (23, 17, 'sp4_v_b_10')
// (23, 17, 'sp4_v_t_47')
// (23, 18, 'sp4_v_b_47')
// (23, 19, 'sp4_v_b_34')
// (23, 20, 'sp4_v_b_23')
// (23, 21, 'sp4_v_b_10')
// (23, 21, 'sp4_v_t_43')
// (23, 22, 'local_g3_3')
// (23, 22, 'lutff_global/cen')
// (23, 22, 'sp4_v_b_43')
// (23, 23, 'sp4_v_b_30')
// (23, 24, 'sp4_v_b_19')
// (23, 25, 'sp4_v_b_6')
// (24, 13, 'sp4_h_r_23')
// (25, 13, 'sp4_h_r_34')
// (26, 13, 'sp4_h_r_47')
// (27, 13, 'sp4_h_l_47')

wire n794;
// (14, 14, 'sp4_r_v_b_43')
// (14, 15, 'sp4_r_v_b_30')
// (14, 16, 'sp4_r_v_b_19')
// (14, 17, 'local_g1_6')
// (14, 17, 'lutff_4/in_1')
// (14, 17, 'sp4_r_v_b_6')
// (15, 13, 'sp4_h_r_0')
// (15, 13, 'sp4_v_t_43')
// (15, 14, 'sp4_v_b_43')
// (15, 15, 'sp4_v_b_30')
// (15, 16, 'sp4_v_b_19')
// (15, 17, 'sp4_v_b_6')
// (16, 12, 'neigh_op_tnr_4')
// (16, 13, 'neigh_op_rgt_4')
// (16, 13, 'sp4_h_r_13')
// (16, 14, 'neigh_op_bnr_4')
// (17, 12, 'neigh_op_top_4')
// (17, 13, 'lutff_4/out')
// (17, 13, 'sp4_h_r_24')
// (17, 14, 'neigh_op_bot_4')
// (18, 12, 'neigh_op_tnl_4')
// (18, 13, 'neigh_op_lft_4')
// (18, 13, 'sp4_h_r_37')
// (18, 14, 'neigh_op_bnl_4')
// (19, 13, 'sp4_h_l_37')

reg n795 = 0;
// (14, 14, 'sp4_r_v_b_45')
// (14, 15, 'sp4_r_v_b_32')
// (14, 16, 'sp4_r_v_b_21')
// (14, 17, 'local_g2_0')
// (14, 17, 'lutff_5/in_1')
// (14, 17, 'sp4_r_v_b_8')
// (15, 13, 'sp4_h_r_8')
// (15, 13, 'sp4_v_t_45')
// (15, 14, 'sp4_v_b_45')
// (15, 15, 'sp4_v_b_32')
// (15, 16, 'sp4_v_b_21')
// (15, 17, 'sp4_v_b_8')
// (16, 13, 'sp4_h_r_21')
// (17, 13, 'sp4_h_r_32')
// (18, 13, 'sp4_h_r_45')
// (19, 13, 'sp4_h_l_45')
// (19, 13, 'sp4_h_r_8')
// (20, 13, 'sp4_h_r_21')
// (21, 13, 'sp4_h_r_32')
// (22, 10, 'sp4_r_v_b_38')
// (22, 11, 'neigh_op_tnr_7')
// (22, 11, 'sp4_r_v_b_27')
// (22, 12, 'neigh_op_rgt_7')
// (22, 12, 'sp4_r_v_b_14')
// (22, 13, 'neigh_op_bnr_7')
// (22, 13, 'sp4_h_r_45')
// (22, 13, 'sp4_r_v_b_3')
// (23, 9, 'sp4_v_t_38')
// (23, 10, 'sp4_v_b_38')
// (23, 11, 'neigh_op_top_7')
// (23, 11, 'sp4_v_b_27')
// (23, 12, 'lutff_7/out')
// (23, 12, 'sp4_v_b_14')
// (23, 13, 'neigh_op_bot_7')
// (23, 13, 'sp4_h_l_45')
// (23, 13, 'sp4_v_b_3')
// (24, 11, 'neigh_op_tnl_7')
// (24, 12, 'neigh_op_lft_7')
// (24, 13, 'neigh_op_bnl_7')

reg n796 = 0;
// (14, 15, 'local_g2_5')
// (14, 15, 'lutff_0/in_3')
// (14, 15, 'sp4_r_v_b_37')
// (14, 16, 'sp4_r_v_b_24')
// (14, 17, 'sp4_r_v_b_13')
// (14, 18, 'sp4_r_v_b_0')
// (14, 19, 'sp4_r_v_b_41')
// (14, 20, 'sp4_r_v_b_28')
// (14, 21, 'sp4_r_v_b_17')
// (14, 22, 'sp4_r_v_b_4')
// (15, 14, 'sp4_v_t_37')
// (15, 15, 'sp4_v_b_37')
// (15, 16, 'sp4_v_b_24')
// (15, 17, 'sp4_v_b_13')
// (15, 18, 'sp4_v_b_0')
// (15, 18, 'sp4_v_t_41')
// (15, 19, 'sp4_v_b_41')
// (15, 20, 'sp4_v_b_28')
// (15, 21, 'sp4_v_b_17')
// (15, 22, 'sp4_h_r_4')
// (15, 22, 'sp4_v_b_4')
// (16, 22, 'sp4_h_r_17')
// (17, 22, 'sp4_h_r_28')
// (18, 22, 'sp4_h_r_41')
// (18, 23, 'neigh_op_tnr_6')
// (18, 23, 'sp4_r_v_b_41')
// (18, 24, 'neigh_op_rgt_6')
// (18, 24, 'sp4_r_v_b_28')
// (18, 25, 'neigh_op_bnr_6')
// (18, 25, 'sp4_r_v_b_17')
// (18, 26, 'sp4_r_v_b_4')
// (19, 22, 'sp4_h_l_41')
// (19, 22, 'sp4_v_t_41')
// (19, 23, 'neigh_op_top_6')
// (19, 23, 'sp4_v_b_41')
// (19, 24, 'local_g1_6')
// (19, 24, 'lutff_6/in_1')
// (19, 24, 'lutff_6/out')
// (19, 24, 'sp4_v_b_28')
// (19, 25, 'neigh_op_bot_6')
// (19, 25, 'sp4_v_b_17')
// (19, 26, 'sp4_v_b_4')
// (20, 23, 'neigh_op_tnl_6')
// (20, 24, 'neigh_op_lft_6')
// (20, 25, 'neigh_op_bnl_6')

reg n797 = 0;
// (14, 15, 'local_g2_7')
// (14, 15, 'lutff_0/in_1')
// (14, 15, 'sp4_r_v_b_39')
// (14, 16, 'sp4_r_v_b_26')
// (14, 17, 'sp4_r_v_b_15')
// (14, 18, 'sp4_r_v_b_2')
// (14, 19, 'sp4_r_v_b_43')
// (14, 20, 'sp4_r_v_b_30')
// (14, 21, 'sp4_r_v_b_19')
// (14, 22, 'sp4_r_v_b_6')
// (15, 14, 'sp4_v_t_39')
// (15, 15, 'sp4_v_b_39')
// (15, 16, 'sp4_v_b_26')
// (15, 17, 'sp4_v_b_15')
// (15, 18, 'sp4_v_b_2')
// (15, 18, 'sp4_v_t_43')
// (15, 19, 'sp4_v_b_43')
// (15, 20, 'sp4_v_b_30')
// (15, 21, 'sp4_v_b_19')
// (15, 22, 'sp4_h_r_6')
// (15, 22, 'sp4_v_b_6')
// (16, 22, 'sp4_h_r_19')
// (17, 22, 'sp4_h_r_30')
// (18, 22, 'sp4_h_r_43')
// (18, 23, 'neigh_op_tnr_7')
// (18, 23, 'sp4_r_v_b_43')
// (18, 24, 'neigh_op_rgt_7')
// (18, 24, 'sp4_r_v_b_30')
// (18, 25, 'neigh_op_bnr_7')
// (18, 25, 'sp4_r_v_b_19')
// (18, 26, 'sp4_r_v_b_6')
// (19, 22, 'sp4_h_l_43')
// (19, 22, 'sp4_v_t_43')
// (19, 23, 'neigh_op_top_7')
// (19, 23, 'sp4_v_b_43')
// (19, 24, 'local_g1_7')
// (19, 24, 'lutff_7/in_1')
// (19, 24, 'lutff_7/out')
// (19, 24, 'sp4_v_b_30')
// (19, 25, 'neigh_op_bot_7')
// (19, 25, 'sp4_v_b_19')
// (19, 26, 'sp4_v_b_6')
// (20, 23, 'neigh_op_tnl_7')
// (20, 24, 'neigh_op_lft_7')
// (20, 25, 'neigh_op_bnl_7')

wire n798;
// (14, 15, 'lutff_5/lout')
// (14, 15, 'lutff_6/in_2')

wire n799;
// (14, 15, 'neigh_op_tnr_2')
// (14, 16, 'neigh_op_rgt_2')
// (14, 17, 'neigh_op_bnr_2')
// (15, 15, 'neigh_op_top_2')
// (15, 16, 'lutff_2/out')
// (15, 17, 'neigh_op_bot_2')
// (16, 15, 'neigh_op_tnl_2')
// (16, 16, 'local_g0_2')
// (16, 16, 'lutff_global/cen')
// (16, 16, 'neigh_op_lft_2')
// (16, 17, 'neigh_op_bnl_2')

wire n800;
// (14, 15, 'neigh_op_tnr_5')
// (14, 16, 'neigh_op_rgt_5')
// (14, 17, 'neigh_op_bnr_5')
// (15, 15, 'neigh_op_top_5')
// (15, 16, 'lutff_5/out')
// (15, 16, 'sp4_r_v_b_43')
// (15, 17, 'neigh_op_bot_5')
// (15, 17, 'sp4_r_v_b_30')
// (15, 18, 'sp4_r_v_b_19')
// (15, 19, 'sp4_r_v_b_6')
// (16, 15, 'neigh_op_tnl_5')
// (16, 15, 'sp4_v_t_43')
// (16, 16, 'neigh_op_lft_5')
// (16, 16, 'sp4_v_b_43')
// (16, 17, 'neigh_op_bnl_5')
// (16, 17, 'sp4_v_b_30')
// (16, 18, 'local_g1_3')
// (16, 18, 'lutff_global/cen')
// (16, 18, 'sp4_v_b_19')
// (16, 19, 'sp4_v_b_6')

wire n801;
// (14, 15, 'neigh_op_tnr_7')
// (14, 16, 'neigh_op_rgt_7')
// (14, 17, 'neigh_op_bnr_7')
// (15, 15, 'neigh_op_top_7')
// (15, 15, 'sp4_r_v_b_42')
// (15, 16, 'lutff_7/out')
// (15, 16, 'sp4_r_v_b_31')
// (15, 17, 'neigh_op_bot_7')
// (15, 17, 'sp4_r_v_b_18')
// (15, 18, 'sp4_r_v_b_7')
// (15, 19, 'sp4_r_v_b_42')
// (15, 20, 'sp4_r_v_b_31')
// (15, 21, 'sp4_r_v_b_18')
// (15, 22, 'sp4_r_v_b_7')
// (16, 14, 'sp4_v_t_42')
// (16, 15, 'neigh_op_tnl_7')
// (16, 15, 'sp4_v_b_42')
// (16, 16, 'neigh_op_lft_7')
// (16, 16, 'sp4_v_b_31')
// (16, 17, 'neigh_op_bnl_7')
// (16, 17, 'sp4_v_b_18')
// (16, 18, 'sp4_v_b_7')
// (16, 18, 'sp4_v_t_42')
// (16, 19, 'local_g2_2')
// (16, 19, 'lutff_global/cen')
// (16, 19, 'sp4_v_b_42')
// (16, 20, 'sp4_v_b_31')
// (16, 21, 'sp4_v_b_18')
// (16, 22, 'sp4_v_b_7')

wire n802;
// (14, 15, 'sp12_h_r_0')
// (15, 14, 'neigh_op_tnr_6')
// (15, 15, 'neigh_op_rgt_6')
// (15, 15, 'sp12_h_r_3')
// (15, 16, 'neigh_op_bnr_6')
// (16, 13, 'sp4_r_v_b_37')
// (16, 14, 'neigh_op_top_6')
// (16, 14, 'sp4_r_v_b_24')
// (16, 15, 'local_g2_6')
// (16, 15, 'lutff_1/in_1')
// (16, 15, 'lutff_2/in_2')
// (16, 15, 'lutff_4/in_0')
// (16, 15, 'lutff_6/out')
// (16, 15, 'sp12_h_r_4')
// (16, 15, 'sp4_r_v_b_13')
// (16, 16, 'neigh_op_bot_6')
// (16, 16, 'sp4_r_v_b_0')
// (17, 12, 'sp4_h_r_0')
// (17, 12, 'sp4_v_t_37')
// (17, 13, 'sp4_v_b_37')
// (17, 14, 'neigh_op_tnl_6')
// (17, 14, 'sp4_v_b_24')
// (17, 15, 'neigh_op_lft_6')
// (17, 15, 'sp12_h_r_7')
// (17, 15, 'sp4_v_b_13')
// (17, 16, 'neigh_op_bnl_6')
// (17, 16, 'sp4_v_b_0')
// (18, 12, 'sp4_h_r_13')
// (18, 15, 'sp12_h_r_8')
// (19, 12, 'local_g2_0')
// (19, 12, 'local_g3_0')
// (19, 12, 'lutff_0/in_2')
// (19, 12, 'lutff_2/in_3')
// (19, 12, 'lutff_3/in_2')
// (19, 12, 'lutff_4/in_0')
// (19, 12, 'sp4_h_r_24')
// (19, 15, 'sp12_h_r_11')
// (20, 12, 'sp4_h_r_37')
// (20, 15, 'sp12_h_r_12')
// (21, 12, 'sp4_h_l_37')
// (21, 15, 'sp12_h_r_15')
// (22, 15, 'local_g0_0')
// (22, 15, 'local_g1_0')
// (22, 15, 'lutff_1/in_2')
// (22, 15, 'lutff_2/in_2')
// (22, 15, 'lutff_3/in_2')
// (22, 15, 'lutff_4/in_2')
// (22, 15, 'sp12_h_r_16')
// (23, 15, 'sp12_h_r_19')
// (24, 15, 'sp12_h_r_20')
// (25, 15, 'sp12_h_r_23')
// (26, 15, 'sp12_h_l_23')

wire n803;
// (14, 15, 'sp4_h_r_0')
// (15, 14, 'neigh_op_tnr_4')
// (15, 15, 'neigh_op_rgt_4')
// (15, 15, 'sp4_h_r_13')
// (15, 16, 'neigh_op_bnr_4')
// (16, 14, 'neigh_op_top_4')
// (16, 15, 'lutff_4/out')
// (16, 15, 'sp4_h_r_24')
// (16, 16, 'neigh_op_bot_4')
// (17, 14, 'neigh_op_tnl_4')
// (17, 15, 'neigh_op_lft_4')
// (17, 15, 'sp4_h_r_37')
// (17, 16, 'neigh_op_bnl_4')
// (17, 16, 'sp4_r_v_b_40')
// (17, 17, 'sp4_r_v_b_29')
// (17, 18, 'sp4_r_v_b_16')
// (17, 19, 'sp4_r_v_b_5')
// (18, 15, 'sp4_h_l_37')
// (18, 15, 'sp4_v_t_40')
// (18, 16, 'sp4_v_b_40')
// (18, 17, 'sp4_v_b_29')
// (18, 18, 'sp4_v_b_16')
// (18, 19, 'sp4_h_r_11')
// (18, 19, 'sp4_v_b_5')
// (19, 19, 'sp4_h_r_22')
// (20, 19, 'local_g3_3')
// (20, 19, 'lutff_global/cen')
// (20, 19, 'sp4_h_r_35')
// (21, 19, 'sp4_h_r_46')
// (22, 19, 'sp4_h_l_46')

reg n804 = 0;
// (14, 15, 'sp4_h_r_5')
// (15, 15, 'sp4_h_r_16')
// (16, 15, 'sp4_h_r_29')
// (17, 15, 'local_g3_0')
// (17, 15, 'lutff_0/in_1')
// (17, 15, 'sp4_h_r_40')
// (18, 15, 'sp4_h_l_40')
// (18, 15, 'sp4_h_r_9')
// (19, 15, 'sp4_h_r_20')
// (20, 15, 'sp4_h_r_33')
// (21, 11, 'neigh_op_tnr_6')
// (21, 12, 'neigh_op_rgt_6')
// (21, 12, 'sp4_r_v_b_44')
// (21, 13, 'neigh_op_bnr_6')
// (21, 13, 'sp4_r_v_b_33')
// (21, 14, 'sp4_r_v_b_20')
// (21, 15, 'sp4_h_r_44')
// (21, 15, 'sp4_r_v_b_9')
// (22, 11, 'neigh_op_top_6')
// (22, 11, 'sp4_v_t_44')
// (22, 12, 'lutff_6/out')
// (22, 12, 'sp4_v_b_44')
// (22, 13, 'neigh_op_bot_6')
// (22, 13, 'sp4_v_b_33')
// (22, 14, 'sp4_v_b_20')
// (22, 15, 'sp4_h_l_44')
// (22, 15, 'sp4_v_b_9')
// (23, 11, 'neigh_op_tnl_6')
// (23, 12, 'neigh_op_lft_6')
// (23, 13, 'neigh_op_bnl_6')

wire n805;
// (14, 15, 'sp4_h_r_7')
// (15, 15, 'sp4_h_r_18')
// (16, 14, 'sp4_h_r_3')
// (16, 15, 'sp4_h_r_31')
// (17, 14, 'sp4_h_r_14')
// (17, 15, 'local_g2_2')
// (17, 15, 'lutff_global/cen')
// (17, 15, 'sp4_h_r_42')
// (18, 14, 'sp4_h_r_27')
// (18, 15, 'sp4_h_l_42')
// (18, 15, 'sp4_h_r_4')
// (19, 14, 'neigh_op_tnr_6')
// (19, 14, 'sp4_h_r_38')
// (19, 15, 'neigh_op_rgt_6')
// (19, 15, 'sp4_h_r_17')
// (19, 15, 'sp4_r_v_b_44')
// (19, 16, 'neigh_op_bnr_6')
// (19, 16, 'sp4_r_v_b_33')
// (19, 17, 'sp4_r_v_b_20')
// (19, 18, 'sp4_r_v_b_9')
// (20, 14, 'neigh_op_top_6')
// (20, 14, 'sp4_h_l_38')
// (20, 14, 'sp4_h_r_6')
// (20, 14, 'sp4_v_t_44')
// (20, 15, 'lutff_6/out')
// (20, 15, 'sp4_h_r_28')
// (20, 15, 'sp4_v_b_44')
// (20, 16, 'neigh_op_bot_6')
// (20, 16, 'sp4_v_b_33')
// (20, 17, 'sp4_v_b_20')
// (20, 18, 'sp4_v_b_9')
// (21, 12, 'sp4_r_v_b_47')
// (21, 13, 'sp4_r_v_b_34')
// (21, 14, 'local_g1_3')
// (21, 14, 'lutff_global/cen')
// (21, 14, 'neigh_op_tnl_6')
// (21, 14, 'sp4_h_r_19')
// (21, 14, 'sp4_r_v_b_23')
// (21, 15, 'neigh_op_lft_6')
// (21, 15, 'sp4_h_r_41')
// (21, 15, 'sp4_r_v_b_10')
// (21, 16, 'neigh_op_bnl_6')
// (22, 11, 'sp4_v_t_47')
// (22, 12, 'sp4_v_b_47')
// (22, 13, 'local_g2_2')
// (22, 13, 'lutff_global/cen')
// (22, 13, 'sp4_v_b_34')
// (22, 14, 'sp4_h_r_30')
// (22, 14, 'sp4_v_b_23')
// (22, 15, 'sp4_h_l_41')
// (22, 15, 'sp4_v_b_10')
// (23, 11, 'sp4_r_v_b_43')
// (23, 12, 'sp4_r_v_b_30')
// (23, 13, 'sp4_r_v_b_19')
// (23, 14, 'sp4_h_r_43')
// (23, 14, 'sp4_r_v_b_6')
// (24, 10, 'sp4_v_t_43')
// (24, 11, 'sp4_v_b_43')
// (24, 12, 'sp4_v_b_30')
// (24, 13, 'local_g1_3')
// (24, 13, 'lutff_global/cen')
// (24, 13, 'sp4_v_b_19')
// (24, 14, 'sp4_h_l_43')
// (24, 14, 'sp4_v_b_6')

reg n806 = 0;
// (14, 15, 'sp4_r_v_b_36')
// (14, 16, 'neigh_op_tnr_6')
// (14, 16, 'sp4_r_v_b_25')
// (14, 17, 'neigh_op_rgt_6')
// (14, 17, 'sp4_r_v_b_12')
// (14, 18, 'neigh_op_bnr_6')
// (14, 18, 'sp4_r_v_b_1')
// (15, 14, 'sp4_h_r_1')
// (15, 14, 'sp4_v_t_36')
// (15, 15, 'sp4_v_b_36')
// (15, 16, 'neigh_op_top_6')
// (15, 16, 'sp4_v_b_25')
// (15, 17, 'lutff_6/out')
// (15, 17, 'sp4_v_b_12')
// (15, 18, 'neigh_op_bot_6')
// (15, 18, 'sp4_v_b_1')
// (16, 14, 'sp4_h_r_12')
// (16, 16, 'neigh_op_tnl_6')
// (16, 17, 'neigh_op_lft_6')
// (16, 18, 'neigh_op_bnl_6')
// (17, 14, 'local_g2_1')
// (17, 14, 'lutff_4/in_1')
// (17, 14, 'sp4_h_r_25')
// (18, 14, 'sp4_h_r_36')
// (19, 14, 'sp4_h_l_36')

wire n807;
// (14, 16, 'lutff_4/lout')
// (14, 16, 'lutff_5/in_2')

reg n808 = 0;
// (14, 16, 'neigh_op_tnr_0')
// (14, 16, 'sp4_r_v_b_45')
// (14, 17, 'neigh_op_rgt_0')
// (14, 17, 'sp4_r_v_b_32')
// (14, 18, 'neigh_op_bnr_0')
// (14, 18, 'sp4_r_v_b_21')
// (14, 19, 'sp4_r_v_b_8')
// (15, 15, 'sp4_h_r_1')
// (15, 15, 'sp4_v_t_45')
// (15, 16, 'neigh_op_top_0')
// (15, 16, 'sp4_v_b_45')
// (15, 17, 'lutff_0/out')
// (15, 17, 'sp4_v_b_32')
// (15, 18, 'neigh_op_bot_0')
// (15, 18, 'sp4_v_b_21')
// (15, 19, 'sp4_v_b_8')
// (16, 15, 'sp4_h_r_12')
// (16, 16, 'neigh_op_tnl_0')
// (16, 17, 'neigh_op_lft_0')
// (16, 18, 'neigh_op_bnl_0')
// (17, 15, 'local_g2_1')
// (17, 15, 'lutff_6/in_1')
// (17, 15, 'sp4_h_r_25')
// (18, 15, 'sp4_h_r_36')
// (19, 15, 'sp4_h_l_36')

reg n809 = 0;
// (14, 16, 'neigh_op_tnr_1')
// (14, 17, 'neigh_op_rgt_1')
// (14, 17, 'sp4_h_r_7')
// (14, 18, 'neigh_op_bnr_1')
// (15, 16, 'neigh_op_top_1')
// (15, 17, 'lutff_1/out')
// (15, 17, 'sp4_h_r_18')
// (15, 18, 'neigh_op_bot_1')
// (16, 16, 'neigh_op_tnl_1')
// (16, 17, 'neigh_op_lft_1')
// (16, 17, 'sp4_h_r_31')
// (16, 18, 'neigh_op_bnl_1')
// (17, 17, 'local_g2_2')
// (17, 17, 'lutff_0/in_0')
// (17, 17, 'sp4_h_r_42')
// (18, 17, 'sp4_h_l_42')

reg n810 = 0;
// (14, 16, 'neigh_op_tnr_2')
// (14, 17, 'neigh_op_rgt_2')
// (14, 18, 'neigh_op_bnr_2')
// (15, 15, 'sp4_r_v_b_45')
// (15, 16, 'neigh_op_top_2')
// (15, 16, 'sp4_r_v_b_32')
// (15, 17, 'lutff_2/out')
// (15, 17, 'sp4_r_v_b_21')
// (15, 18, 'neigh_op_bot_2')
// (15, 18, 'sp4_r_v_b_8')
// (16, 14, 'sp4_v_t_45')
// (16, 15, 'sp4_v_b_45')
// (16, 16, 'neigh_op_tnl_2')
// (16, 16, 'sp4_v_b_32')
// (16, 17, 'neigh_op_lft_2')
// (16, 17, 'sp4_v_b_21')
// (16, 18, 'neigh_op_bnl_2')
// (16, 18, 'sp4_h_r_2')
// (16, 18, 'sp4_v_b_8')
// (17, 18, 'sp4_h_r_15')
// (18, 18, 'sp4_h_r_26')
// (19, 18, 'sp4_h_r_39')
// (20, 18, 'sp4_h_l_39')
// (20, 18, 'sp4_h_r_10')
// (21, 18, 'local_g1_7')
// (21, 18, 'lutff_1/in_1')
// (21, 18, 'sp4_h_r_23')
// (22, 18, 'sp4_h_r_34')
// (23, 18, 'sp4_h_r_47')
// (24, 18, 'sp4_h_l_47')

reg n811 = 0;
// (14, 16, 'neigh_op_tnr_3')
// (14, 17, 'neigh_op_rgt_3')
// (14, 17, 'sp4_h_r_11')
// (14, 18, 'neigh_op_bnr_3')
// (15, 16, 'neigh_op_top_3')
// (15, 17, 'lutff_3/out')
// (15, 17, 'sp4_h_r_22')
// (15, 18, 'neigh_op_bot_3')
// (16, 16, 'neigh_op_tnl_3')
// (16, 17, 'neigh_op_lft_3')
// (16, 17, 'sp4_h_r_35')
// (16, 18, 'neigh_op_bnl_3')
// (17, 17, 'sp4_h_r_46')
// (18, 17, 'sp4_h_l_46')
// (18, 17, 'sp4_h_r_11')
// (19, 17, 'sp4_h_r_22')
// (20, 17, 'sp4_h_r_35')
// (21, 17, 'sp4_h_r_46')
// (21, 18, 'local_g3_6')
// (21, 18, 'lutff_4/in_1')
// (21, 18, 'sp4_r_v_b_46')
// (21, 19, 'sp4_r_v_b_35')
// (21, 20, 'sp4_r_v_b_22')
// (21, 21, 'sp4_r_v_b_11')
// (22, 17, 'sp4_h_l_46')
// (22, 17, 'sp4_v_t_46')
// (22, 18, 'sp4_v_b_46')
// (22, 19, 'sp4_v_b_35')
// (22, 20, 'sp4_v_b_22')
// (22, 21, 'sp4_v_b_11')

reg n812 = 0;
// (14, 16, 'neigh_op_tnr_4')
// (14, 17, 'neigh_op_rgt_4')
// (14, 18, 'neigh_op_bnr_4')
// (15, 16, 'neigh_op_top_4')
// (15, 17, 'lutff_4/out')
// (15, 17, 'sp12_h_r_0')
// (15, 18, 'neigh_op_bot_4')
// (16, 16, 'neigh_op_tnl_4')
// (16, 17, 'neigh_op_lft_4')
// (16, 17, 'sp12_h_r_3')
// (16, 18, 'neigh_op_bnl_4')
// (17, 17, 'sp12_h_r_4')
// (18, 17, 'sp12_h_r_7')
// (19, 17, 'sp12_h_r_8')
// (20, 17, 'sp12_h_r_11')
// (21, 17, 'sp12_h_r_12')
// (21, 18, 'local_g3_4')
// (21, 18, 'lutff_7/in_0')
// (21, 18, 'sp4_r_v_b_44')
// (21, 19, 'sp4_r_v_b_33')
// (21, 20, 'sp4_r_v_b_20')
// (21, 21, 'sp4_r_v_b_9')
// (22, 17, 'sp12_h_r_15')
// (22, 17, 'sp4_h_r_9')
// (22, 17, 'sp4_v_t_44')
// (22, 18, 'sp4_v_b_44')
// (22, 19, 'sp4_v_b_33')
// (22, 20, 'sp4_v_b_20')
// (22, 21, 'sp4_v_b_9')
// (23, 17, 'sp12_h_r_16')
// (23, 17, 'sp4_h_r_20')
// (24, 17, 'sp12_h_r_19')
// (24, 17, 'sp4_h_r_33')
// (25, 17, 'sp12_h_r_20')
// (25, 17, 'sp4_h_r_44')
// (26, 17, 'sp12_h_r_23')
// (26, 17, 'sp4_h_l_44')
// (27, 17, 'sp12_h_l_23')

reg n813 = 0;
// (14, 16, 'neigh_op_tnr_7')
// (14, 17, 'neigh_op_rgt_7')
// (14, 18, 'neigh_op_bnr_7')
// (15, 16, 'neigh_op_top_7')
// (15, 16, 'sp4_r_v_b_42')
// (15, 17, 'lutff_7/out')
// (15, 17, 'sp4_r_v_b_31')
// (15, 18, 'neigh_op_bot_7')
// (15, 18, 'sp4_r_v_b_18')
// (15, 19, 'sp4_r_v_b_7')
// (16, 15, 'sp4_h_r_0')
// (16, 15, 'sp4_v_t_42')
// (16, 16, 'neigh_op_tnl_7')
// (16, 16, 'sp4_v_b_42')
// (16, 17, 'neigh_op_lft_7')
// (16, 17, 'sp4_v_b_31')
// (16, 18, 'neigh_op_bnl_7')
// (16, 18, 'sp4_v_b_18')
// (16, 19, 'sp4_v_b_7')
// (17, 15, 'local_g0_5')
// (17, 15, 'lutff_4/in_3')
// (17, 15, 'sp4_h_r_13')
// (18, 15, 'sp4_h_r_24')
// (19, 15, 'sp4_h_r_37')
// (20, 15, 'sp4_h_l_37')

reg n814 = 0;
// (14, 16, 'sp4_h_r_8')
// (15, 15, 'neigh_op_tnr_0')
// (15, 16, 'neigh_op_rgt_0')
// (15, 16, 'sp4_h_r_21')
// (15, 17, 'neigh_op_bnr_0')
// (16, 15, 'neigh_op_top_0')
// (16, 16, 'lutff_0/out')
// (16, 16, 'sp4_h_r_32')
// (16, 17, 'neigh_op_bot_0')
// (17, 13, 'sp4_r_v_b_45')
// (17, 14, 'sp4_r_v_b_32')
// (17, 15, 'neigh_op_tnl_0')
// (17, 15, 'sp4_r_v_b_21')
// (17, 16, 'neigh_op_lft_0')
// (17, 16, 'sp4_h_r_45')
// (17, 16, 'sp4_r_v_b_8')
// (17, 17, 'neigh_op_bnl_0')
// (18, 12, 'sp4_v_t_45')
// (18, 13, 'sp4_v_b_45')
// (18, 14, 'sp4_v_b_32')
// (18, 15, 'local_g1_5')
// (18, 15, 'lutff_3/in_3')
// (18, 15, 'sp4_v_b_21')
// (18, 16, 'sp4_h_l_45')
// (18, 16, 'sp4_v_b_8')

reg n815 = 0;
// (14, 16, 'sp4_r_v_b_40')
// (14, 17, 'neigh_op_tnr_0')
// (14, 17, 'sp4_r_v_b_29')
// (14, 18, 'neigh_op_rgt_0')
// (14, 18, 'sp4_r_v_b_16')
// (14, 19, 'neigh_op_bnr_0')
// (14, 19, 'sp4_r_v_b_5')
// (15, 15, 'sp4_v_t_40')
// (15, 16, 'sp4_v_b_40')
// (15, 17, 'neigh_op_top_0')
// (15, 17, 'sp4_v_b_29')
// (15, 18, 'lutff_0/out')
// (15, 18, 'sp4_v_b_16')
// (15, 19, 'neigh_op_bot_0')
// (15, 19, 'sp4_h_r_11')
// (15, 19, 'sp4_v_b_5')
// (16, 17, 'neigh_op_tnl_0')
// (16, 18, 'neigh_op_lft_0')
// (16, 19, 'neigh_op_bnl_0')
// (16, 19, 'sp4_h_r_22')
// (17, 19, 'sp4_h_r_35')
// (18, 19, 'local_g3_6')
// (18, 19, 'lutff_2/in_1')
// (18, 19, 'sp4_h_r_46')
// (19, 19, 'sp4_h_l_46')

wire n816;
// (14, 17, 'local_g3_1')
// (14, 17, 'lutff_3/in_1')
// (14, 17, 'sp4_r_v_b_41')
// (14, 18, 'sp4_r_v_b_28')
// (14, 19, 'sp4_r_v_b_17')
// (14, 20, 'sp4_r_v_b_4')
// (15, 16, 'sp4_v_t_41')
// (15, 17, 'sp4_v_b_41')
// (15, 18, 'sp4_v_b_28')
// (15, 19, 'sp4_v_b_17')
// (15, 20, 'sp4_h_r_11')
// (15, 20, 'sp4_v_b_4')
// (16, 20, 'sp4_h_r_22')
// (17, 20, 'sp4_h_r_35')
// (17, 23, 'neigh_op_tnr_5')
// (17, 24, 'neigh_op_rgt_5')
// (17, 25, 'neigh_op_bnr_5')
// (18, 20, 'sp4_h_r_46')
// (18, 21, 'sp4_r_v_b_46')
// (18, 22, 'sp4_r_v_b_35')
// (18, 23, 'neigh_op_top_5')
// (18, 23, 'sp4_r_v_b_22')
// (18, 24, 'lutff_5/out')
// (18, 24, 'sp4_r_v_b_11')
// (18, 25, 'neigh_op_bot_5')
// (19, 20, 'sp4_h_l_46')
// (19, 20, 'sp4_v_t_46')
// (19, 21, 'sp4_v_b_46')
// (19, 22, 'sp4_v_b_35')
// (19, 23, 'neigh_op_tnl_5')
// (19, 23, 'sp4_v_b_22')
// (19, 24, 'neigh_op_lft_5')
// (19, 24, 'sp4_v_b_11')
// (19, 25, 'neigh_op_bnl_5')

wire n817;
// (14, 17, 'lutff_3/lout')
// (14, 17, 'lutff_4/in_2')

wire n818;
// (14, 17, 'lutff_4/lout')
// (14, 17, 'lutff_5/in_2')

reg n819 = 0;
// (14, 17, 'neigh_op_tnr_2')
// (14, 18, 'neigh_op_rgt_2')
// (14, 19, 'neigh_op_bnr_2')
// (15, 17, 'neigh_op_top_2')
// (15, 18, 'lutff_2/out')
// (15, 18, 'sp4_h_r_4')
// (15, 19, 'neigh_op_bot_2')
// (16, 17, 'neigh_op_tnl_2')
// (16, 18, 'neigh_op_lft_2')
// (16, 18, 'sp4_h_r_17')
// (16, 19, 'neigh_op_bnl_2')
// (17, 18, 'sp4_h_r_28')
// (18, 18, 'sp4_h_r_41')
// (19, 18, 'sp4_h_l_41')
// (19, 18, 'sp4_h_r_0')
// (20, 18, 'sp4_h_r_13')
// (21, 18, 'sp4_h_r_24')
// (22, 18, 'sp4_h_r_37')
// (22, 19, 'sp4_r_v_b_37')
// (22, 20, 'local_g0_0')
// (22, 20, 'lutff_7/in_1')
// (22, 20, 'sp4_r_v_b_24')
// (22, 21, 'sp4_r_v_b_13')
// (22, 22, 'sp4_r_v_b_0')
// (23, 18, 'sp4_h_l_37')
// (23, 18, 'sp4_v_t_37')
// (23, 19, 'sp4_v_b_37')
// (23, 20, 'sp4_v_b_24')
// (23, 21, 'sp4_v_b_13')
// (23, 22, 'sp4_v_b_0')

reg n820 = 0;
// (14, 17, 'neigh_op_tnr_3')
// (14, 18, 'neigh_op_rgt_3')
// (14, 19, 'neigh_op_bnr_3')
// (15, 16, 'sp4_r_v_b_47')
// (15, 17, 'neigh_op_top_3')
// (15, 17, 'sp4_r_v_b_34')
// (15, 18, 'lutff_3/out')
// (15, 18, 'sp4_r_v_b_23')
// (15, 19, 'neigh_op_bot_3')
// (15, 19, 'sp4_r_v_b_10')
// (16, 15, 'sp4_v_t_47')
// (16, 16, 'sp4_v_b_47')
// (16, 17, 'neigh_op_tnl_3')
// (16, 17, 'sp4_v_b_34')
// (16, 18, 'neigh_op_lft_3')
// (16, 18, 'sp4_v_b_23')
// (16, 19, 'neigh_op_bnl_3')
// (16, 19, 'sp4_h_r_10')
// (16, 19, 'sp4_v_b_10')
// (17, 19, 'sp4_h_r_23')
// (18, 19, 'local_g2_2')
// (18, 19, 'lutff_3/in_1')
// (18, 19, 'sp4_h_r_34')
// (19, 19, 'sp4_h_r_47')
// (20, 19, 'sp4_h_l_47')

reg n821 = 0;
// (14, 17, 'neigh_op_tnr_4')
// (14, 18, 'neigh_op_rgt_4')
// (14, 19, 'neigh_op_bnr_4')
// (15, 17, 'neigh_op_top_4')
// (15, 17, 'sp4_r_v_b_36')
// (15, 18, 'lutff_4/out')
// (15, 18, 'sp4_r_v_b_25')
// (15, 19, 'neigh_op_bot_4')
// (15, 19, 'sp4_r_v_b_12')
// (15, 20, 'sp4_r_v_b_1')
// (16, 16, 'sp4_v_t_36')
// (16, 17, 'neigh_op_tnl_4')
// (16, 17, 'sp4_v_b_36')
// (16, 18, 'neigh_op_lft_4')
// (16, 18, 'sp4_v_b_25')
// (16, 19, 'neigh_op_bnl_4')
// (16, 19, 'sp4_v_b_12')
// (16, 20, 'sp4_h_r_1')
// (16, 20, 'sp4_v_b_1')
// (17, 20, 'sp4_h_r_12')
// (18, 20, 'local_g3_1')
// (18, 20, 'lutff_5/in_1')
// (18, 20, 'sp4_h_r_25')
// (19, 20, 'sp4_h_r_36')
// (20, 20, 'sp4_h_l_36')

reg n822 = 0;
// (14, 17, 'neigh_op_tnr_5')
// (14, 18, 'neigh_op_rgt_5')
// (14, 19, 'neigh_op_bnr_5')
// (15, 17, 'neigh_op_top_5')
// (15, 18, 'lutff_5/out')
// (15, 18, 'sp4_h_r_10')
// (15, 19, 'neigh_op_bot_5')
// (16, 17, 'neigh_op_tnl_5')
// (16, 18, 'neigh_op_lft_5')
// (16, 18, 'sp4_h_r_23')
// (16, 19, 'neigh_op_bnl_5')
// (17, 18, 'sp4_h_r_34')
// (18, 18, 'local_g3_7')
// (18, 18, 'lutff_0/in_0')
// (18, 18, 'sp4_h_r_47')
// (19, 18, 'sp4_h_l_47')

reg n823 = 0;
// (14, 17, 'neigh_op_tnr_6')
// (14, 18, 'neigh_op_rgt_6')
// (14, 19, 'neigh_op_bnr_6')
// (15, 16, 'sp4_r_v_b_37')
// (15, 17, 'neigh_op_top_6')
// (15, 17, 'sp4_r_v_b_24')
// (15, 18, 'lutff_6/out')
// (15, 18, 'sp4_r_v_b_13')
// (15, 19, 'neigh_op_bot_6')
// (15, 19, 'sp4_r_v_b_0')
// (16, 15, 'sp4_v_t_37')
// (16, 16, 'sp4_v_b_37')
// (16, 17, 'neigh_op_tnl_6')
// (16, 17, 'sp4_v_b_24')
// (16, 18, 'neigh_op_lft_6')
// (16, 18, 'sp4_v_b_13')
// (16, 19, 'neigh_op_bnl_6')
// (16, 19, 'sp4_h_r_0')
// (16, 19, 'sp4_v_b_0')
// (17, 19, 'sp4_h_r_13')
// (18, 19, 'local_g3_0')
// (18, 19, 'lutff_4/in_1')
// (18, 19, 'sp4_h_r_24')
// (19, 19, 'sp4_h_r_37')
// (20, 19, 'sp4_h_l_37')

reg n824 = 0;
// (14, 17, 'neigh_op_tnr_7')
// (14, 18, 'neigh_op_rgt_7')
// (14, 19, 'neigh_op_bnr_7')
// (15, 17, 'neigh_op_top_7')
// (15, 18, 'lutff_7/out')
// (15, 18, 'sp4_r_v_b_47')
// (15, 19, 'neigh_op_bot_7')
// (15, 19, 'sp4_r_v_b_34')
// (15, 20, 'sp4_r_v_b_23')
// (15, 21, 'sp4_r_v_b_10')
// (16, 17, 'neigh_op_tnl_7')
// (16, 17, 'sp4_h_r_10')
// (16, 17, 'sp4_v_t_47')
// (16, 18, 'neigh_op_lft_7')
// (16, 18, 'sp4_v_b_47')
// (16, 19, 'neigh_op_bnl_7')
// (16, 19, 'sp4_v_b_34')
// (16, 20, 'sp4_v_b_23')
// (16, 21, 'sp4_v_b_10')
// (17, 17, 'sp4_h_r_23')
// (18, 17, 'local_g2_2')
// (18, 17, 'lutff_0/in_0')
// (18, 17, 'sp4_h_r_34')
// (19, 17, 'sp4_h_r_47')
// (20, 17, 'sp4_h_l_47')

reg n825 = 0;
// (14, 17, 'sp4_h_r_0')
// (15, 16, 'neigh_op_tnr_4')
// (15, 17, 'neigh_op_rgt_4')
// (15, 17, 'sp4_h_r_13')
// (15, 18, 'neigh_op_bnr_4')
// (16, 16, 'neigh_op_top_4')
// (16, 17, 'lutff_4/out')
// (16, 17, 'sp4_h_r_24')
// (16, 18, 'neigh_op_bot_4')
// (17, 16, 'neigh_op_tnl_4')
// (17, 17, 'neigh_op_lft_4')
// (17, 17, 'sp4_h_r_37')
// (17, 18, 'neigh_op_bnl_4')
// (18, 17, 'sp4_h_l_37')
// (18, 17, 'sp4_h_r_0')
// (19, 17, 'sp4_h_r_13')
// (20, 17, 'sp4_h_r_24')
// (21, 17, 'sp4_h_r_37')
// (21, 18, 'local_g3_0')
// (21, 18, 'lutff_6/in_1')
// (21, 18, 'sp4_r_v_b_40')
// (21, 19, 'sp4_r_v_b_29')
// (21, 20, 'sp4_r_v_b_16')
// (21, 21, 'sp4_r_v_b_5')
// (22, 17, 'sp4_h_l_37')
// (22, 17, 'sp4_v_t_40')
// (22, 18, 'sp4_v_b_40')
// (22, 19, 'sp4_v_b_29')
// (22, 20, 'sp4_v_b_16')
// (22, 21, 'sp4_v_b_5')

wire n826;
// (14, 17, 'sp4_r_v_b_39')
// (14, 18, 'sp4_r_v_b_26')
// (14, 19, 'sp4_r_v_b_15')
// (14, 20, 'sp4_r_v_b_2')
// (15, 16, 'sp4_v_t_39')
// (15, 17, 'sp4_v_b_39')
// (15, 18, 'local_g2_2')
// (15, 18, 'lutff_global/cen')
// (15, 18, 'sp4_v_b_26')
// (15, 19, 'neigh_op_tnr_2')
// (15, 19, 'sp4_v_b_15')
// (15, 20, 'neigh_op_rgt_2')
// (15, 20, 'sp4_h_r_9')
// (15, 20, 'sp4_v_b_2')
// (15, 21, 'neigh_op_bnr_2')
// (16, 19, 'neigh_op_top_2')
// (16, 20, 'lutff_2/out')
// (16, 20, 'sp4_h_r_20')
// (16, 21, 'neigh_op_bot_2')
// (17, 19, 'neigh_op_tnl_2')
// (17, 20, 'neigh_op_lft_2')
// (17, 20, 'sp4_h_r_33')
// (17, 21, 'neigh_op_bnl_2')
// (18, 20, 'sp4_h_r_44')
// (19, 20, 'sp4_h_l_44')

wire n827;
// (14, 18, 'carry_in_mux')
// (14, 18, 'lutff_0/in_3')

wire n828;
// (14, 18, 'lutff_0/cout')
// (14, 18, 'lutff_1/in_3')

wire n829;
// (14, 18, 'lutff_1/cout')
// (14, 18, 'lutff_2/in_3')

wire n830;
// (14, 18, 'lutff_2/cout')
// (14, 18, 'lutff_3/in_3')

wire n831;
// (14, 18, 'lutff_3/cout')
// (14, 18, 'lutff_4/in_3')

wire n832;
// (14, 18, 'lutff_4/cout')
// (14, 18, 'lutff_5/in_3')

wire n833;
// (14, 18, 'lutff_5/cout')
// (14, 18, 'lutff_6/in_3')

wire n834;
// (14, 18, 'lutff_6/cout')
// (14, 18, 'lutff_7/in_3')

wire n835;
// (14, 18, 'lutff_7/cout')
// (14, 19, 'carry_in')
// (14, 19, 'carry_in_mux')
// (14, 19, 'lutff_0/in_3')

reg n836 = 0;
// (14, 18, 'neigh_op_tnr_0')
// (14, 19, 'neigh_op_rgt_0')
// (14, 20, 'neigh_op_bnr_0')
// (15, 18, 'neigh_op_top_0')
// (15, 19, 'lutff_0/out')
// (15, 20, 'local_g1_0')
// (15, 20, 'lutff_0/in_3')
// (15, 20, 'neigh_op_bot_0')
// (16, 18, 'neigh_op_tnl_0')
// (16, 19, 'neigh_op_lft_0')
// (16, 20, 'neigh_op_bnl_0')

reg n837 = 0;
// (14, 18, 'neigh_op_tnr_1')
// (14, 19, 'neigh_op_rgt_1')
// (14, 20, 'neigh_op_bnr_1')
// (15, 18, 'neigh_op_top_1')
// (15, 19, 'lutff_1/out')
// (15, 20, 'local_g0_1')
// (15, 20, 'lutff_1/in_0')
// (15, 20, 'neigh_op_bot_1')
// (16, 18, 'neigh_op_tnl_1')
// (16, 19, 'neigh_op_lft_1')
// (16, 20, 'neigh_op_bnl_1')

reg n838 = 0;
// (14, 18, 'neigh_op_tnr_3')
// (14, 19, 'neigh_op_rgt_3')
// (14, 20, 'neigh_op_bnr_3')
// (15, 18, 'neigh_op_top_3')
// (15, 19, 'lutff_3/out')
// (15, 20, 'local_g1_3')
// (15, 20, 'lutff_3/in_3')
// (15, 20, 'neigh_op_bot_3')
// (16, 18, 'neigh_op_tnl_3')
// (16, 19, 'neigh_op_lft_3')
// (16, 20, 'neigh_op_bnl_3')

reg n839 = 0;
// (14, 18, 'neigh_op_tnr_4')
// (14, 19, 'neigh_op_rgt_4')
// (14, 20, 'neigh_op_bnr_4')
// (15, 18, 'neigh_op_top_4')
// (15, 19, 'lutff_4/out')
// (15, 20, 'local_g1_4')
// (15, 20, 'lutff_4/in_3')
// (15, 20, 'neigh_op_bot_4')
// (16, 18, 'neigh_op_tnl_4')
// (16, 19, 'neigh_op_lft_4')
// (16, 20, 'neigh_op_bnl_4')

reg n840 = 0;
// (14, 18, 'neigh_op_tnr_5')
// (14, 19, 'neigh_op_rgt_5')
// (14, 20, 'neigh_op_bnr_5')
// (15, 18, 'neigh_op_top_5')
// (15, 19, 'lutff_5/out')
// (15, 20, 'local_g0_5')
// (15, 20, 'lutff_5/in_0')
// (15, 20, 'neigh_op_bot_5')
// (16, 18, 'neigh_op_tnl_5')
// (16, 19, 'neigh_op_lft_5')
// (16, 20, 'neigh_op_bnl_5')

reg n841 = 0;
// (14, 18, 'neigh_op_tnr_6')
// (14, 19, 'neigh_op_rgt_6')
// (14, 20, 'neigh_op_bnr_6')
// (15, 18, 'neigh_op_top_6')
// (15, 19, 'lutff_6/out')
// (15, 20, 'local_g1_6')
// (15, 20, 'lutff_6/in_3')
// (15, 20, 'neigh_op_bot_6')
// (16, 18, 'neigh_op_tnl_6')
// (16, 19, 'neigh_op_lft_6')
// (16, 20, 'neigh_op_bnl_6')

reg n842 = 0;
// (14, 18, 'neigh_op_tnr_7')
// (14, 19, 'neigh_op_rgt_7')
// (14, 20, 'neigh_op_bnr_7')
// (15, 18, 'neigh_op_top_7')
// (15, 19, 'lutff_7/out')
// (15, 20, 'local_g1_7')
// (15, 20, 'lutff_7/in_3')
// (15, 20, 'neigh_op_bot_7')
// (16, 18, 'neigh_op_tnl_7')
// (16, 19, 'neigh_op_lft_7')
// (16, 20, 'neigh_op_bnl_7')

reg n843 = 0;
// (14, 18, 'sp4_h_r_10')
// (15, 17, 'neigh_op_tnr_1')
// (15, 18, 'neigh_op_rgt_1')
// (15, 18, 'sp4_h_r_23')
// (15, 19, 'neigh_op_bnr_1')
// (16, 17, 'neigh_op_top_1')
// (16, 18, 'lutff_1/out')
// (16, 18, 'sp4_h_r_34')
// (16, 19, 'neigh_op_bot_1')
// (17, 17, 'neigh_op_tnl_1')
// (17, 18, 'local_g0_1')
// (17, 18, 'lutff_1/in_2')
// (17, 18, 'neigh_op_lft_1')
// (17, 18, 'sp4_h_r_47')
// (17, 19, 'neigh_op_bnl_1')
// (17, 19, 'sp4_r_v_b_47')
// (17, 20, 'sp4_r_v_b_34')
// (17, 21, 'sp4_r_v_b_23')
// (17, 22, 'local_g2_2')
// (17, 22, 'lutff_1/in_3')
// (17, 22, 'sp4_r_v_b_10')
// (18, 18, 'sp4_h_l_47')
// (18, 18, 'sp4_v_t_47')
// (18, 19, 'sp4_v_b_47')
// (18, 20, 'sp4_v_b_34')
// (18, 21, 'sp4_v_b_23')
// (18, 22, 'sp4_v_b_10')

reg n844 = 0;
// (14, 18, 'sp4_h_r_2')
// (15, 17, 'neigh_op_tnr_5')
// (15, 18, 'neigh_op_rgt_5')
// (15, 18, 'sp4_h_r_15')
// (15, 19, 'neigh_op_bnr_5')
// (16, 17, 'neigh_op_top_5')
// (16, 18, 'lutff_5/out')
// (16, 18, 'sp4_h_r_26')
// (16, 19, 'neigh_op_bot_5')
// (17, 17, 'neigh_op_tnl_5')
// (17, 18, 'local_g1_5')
// (17, 18, 'lutff_5/in_1')
// (17, 18, 'neigh_op_lft_5')
// (17, 18, 'sp4_h_r_39')
// (17, 19, 'neigh_op_bnl_5')
// (17, 19, 'sp4_r_v_b_42')
// (17, 20, 'sp4_r_v_b_31')
// (17, 21, 'sp4_r_v_b_18')
// (17, 22, 'local_g1_7')
// (17, 22, 'lutff_5/in_3')
// (17, 22, 'sp4_r_v_b_7')
// (18, 18, 'sp4_h_l_39')
// (18, 18, 'sp4_v_t_42')
// (18, 19, 'sp4_v_b_42')
// (18, 20, 'sp4_v_b_31')
// (18, 21, 'sp4_v_b_18')
// (18, 22, 'sp4_v_b_7')

wire n845;
// (14, 19, 'lutff_0/cout')
// (14, 19, 'lutff_1/in_3')

wire n846;
// (14, 19, 'lutff_1/cout')
// (14, 19, 'lutff_2/in_3')

wire n847;
// (14, 19, 'lutff_2/cout')
// (14, 19, 'lutff_3/in_3')

wire n848;
// (14, 19, 'lutff_3/cout')
// (14, 19, 'lutff_4/in_3')

wire n849;
// (14, 19, 'lutff_4/cout')
// (14, 19, 'lutff_5/in_3')

wire n850;
// (14, 19, 'lutff_5/cout')
// (14, 19, 'lutff_6/in_3')

wire n851;
// (14, 19, 'lutff_6/cout')
// (14, 19, 'lutff_7/in_3')

wire n852;
// (14, 19, 'lutff_7/cout')
// (14, 20, 'carry_in')
// (14, 20, 'carry_in_mux')
// (14, 20, 'lutff_0/in_3')

wire n853;
// (14, 19, 'neigh_op_tnr_0')
// (14, 20, 'neigh_op_rgt_0')
// (14, 21, 'neigh_op_bnr_0')
// (15, 19, 'neigh_op_top_0')
// (15, 20, 'local_g3_0')
// (15, 20, 'lutff_0/in_1')
// (15, 20, 'lutff_0/out')
// (15, 21, 'neigh_op_bot_0')
// (16, 19, 'neigh_op_tnl_0')
// (16, 20, 'neigh_op_lft_0')
// (16, 21, 'neigh_op_bnl_0')

wire n854;
// (14, 19, 'neigh_op_tnr_1')
// (14, 20, 'neigh_op_rgt_1')
// (14, 21, 'neigh_op_bnr_1')
// (15, 19, 'neigh_op_top_1')
// (15, 20, 'local_g3_1')
// (15, 20, 'lutff_1/in_1')
// (15, 20, 'lutff_1/out')
// (15, 21, 'neigh_op_bot_1')
// (16, 19, 'neigh_op_tnl_1')
// (16, 20, 'neigh_op_lft_1')
// (16, 21, 'neigh_op_bnl_1')

wire n855;
// (14, 19, 'neigh_op_tnr_2')
// (14, 20, 'neigh_op_rgt_2')
// (14, 21, 'neigh_op_bnr_2')
// (15, 19, 'neigh_op_top_2')
// (15, 20, 'local_g1_2')
// (15, 20, 'lutff_2/in_1')
// (15, 20, 'lutff_2/out')
// (15, 21, 'neigh_op_bot_2')
// (16, 19, 'neigh_op_tnl_2')
// (16, 20, 'neigh_op_lft_2')
// (16, 21, 'neigh_op_bnl_2')

wire n856;
// (14, 19, 'neigh_op_tnr_3')
// (14, 20, 'neigh_op_rgt_3')
// (14, 21, 'neigh_op_bnr_3')
// (15, 19, 'neigh_op_top_3')
// (15, 20, 'local_g3_3')
// (15, 20, 'lutff_3/in_1')
// (15, 20, 'lutff_3/out')
// (15, 21, 'neigh_op_bot_3')
// (16, 19, 'neigh_op_tnl_3')
// (16, 20, 'neigh_op_lft_3')
// (16, 21, 'neigh_op_bnl_3')

wire n857;
// (14, 19, 'neigh_op_tnr_4')
// (14, 20, 'neigh_op_rgt_4')
// (14, 21, 'neigh_op_bnr_4')
// (15, 19, 'neigh_op_top_4')
// (15, 20, 'local_g3_4')
// (15, 20, 'lutff_4/in_1')
// (15, 20, 'lutff_4/out')
// (15, 21, 'neigh_op_bot_4')
// (16, 19, 'neigh_op_tnl_4')
// (16, 20, 'neigh_op_lft_4')
// (16, 21, 'neigh_op_bnl_4')

wire n858;
// (14, 19, 'neigh_op_tnr_5')
// (14, 20, 'neigh_op_rgt_5')
// (14, 21, 'neigh_op_bnr_5')
// (15, 19, 'neigh_op_top_5')
// (15, 20, 'local_g3_5')
// (15, 20, 'lutff_5/in_1')
// (15, 20, 'lutff_5/out')
// (15, 21, 'neigh_op_bot_5')
// (16, 19, 'neigh_op_tnl_5')
// (16, 20, 'neigh_op_lft_5')
// (16, 21, 'neigh_op_bnl_5')

wire n859;
// (14, 19, 'neigh_op_tnr_6')
// (14, 20, 'neigh_op_rgt_6')
// (14, 21, 'neigh_op_bnr_6')
// (15, 19, 'neigh_op_top_6')
// (15, 20, 'local_g2_6')
// (15, 20, 'lutff_6/in_2')
// (15, 20, 'lutff_6/out')
// (15, 21, 'neigh_op_bot_6')
// (16, 19, 'neigh_op_tnl_6')
// (16, 20, 'neigh_op_lft_6')
// (16, 21, 'neigh_op_bnl_6')

wire n860;
// (14, 19, 'neigh_op_tnr_7')
// (14, 20, 'neigh_op_rgt_7')
// (14, 21, 'neigh_op_bnr_7')
// (15, 19, 'neigh_op_top_7')
// (15, 20, 'local_g3_7')
// (15, 20, 'lutff_7/in_1')
// (15, 20, 'lutff_7/out')
// (15, 21, 'neigh_op_bot_7')
// (16, 19, 'neigh_op_tnl_7')
// (16, 20, 'neigh_op_lft_7')
// (16, 21, 'neigh_op_bnl_7')

reg n861 = 0;
// (14, 19, 'sp4_r_v_b_36')
// (14, 20, 'sp4_r_v_b_25')
// (14, 21, 'sp4_r_v_b_12')
// (14, 22, 'sp4_r_v_b_1')
// (15, 17, 'neigh_op_tnr_6')
// (15, 18, 'neigh_op_rgt_6')
// (15, 18, 'sp4_h_r_1')
// (15, 18, 'sp4_v_t_36')
// (15, 19, 'neigh_op_bnr_6')
// (15, 19, 'sp4_v_b_36')
// (15, 20, 'sp4_v_b_25')
// (15, 21, 'sp4_v_b_12')
// (15, 22, 'sp4_h_r_7')
// (15, 22, 'sp4_v_b_1')
// (16, 17, 'neigh_op_top_6')
// (16, 18, 'lutff_6/out')
// (16, 18, 'sp4_h_r_12')
// (16, 19, 'neigh_op_bot_6')
// (16, 22, 'sp4_h_r_18')
// (17, 17, 'neigh_op_tnl_6')
// (17, 18, 'local_g2_1')
// (17, 18, 'lutff_6/in_1')
// (17, 18, 'neigh_op_lft_6')
// (17, 18, 'sp4_h_r_25')
// (17, 19, 'neigh_op_bnl_6')
// (17, 22, 'local_g2_7')
// (17, 22, 'lutff_6/in_3')
// (17, 22, 'sp4_h_r_31')
// (18, 18, 'sp4_h_r_36')
// (18, 22, 'sp4_h_r_42')
// (19, 18, 'sp4_h_l_36')
// (19, 22, 'sp4_h_l_42')

wire n862;
// (14, 20, 'lutff_0/cout')
// (14, 20, 'lutff_1/in_3')

wire n863;
// (14, 20, 'lutff_1/cout')
// (14, 20, 'lutff_2/in_3')

wire n864;
// (14, 20, 'lutff_2/cout')
// (14, 20, 'lutff_3/in_3')

wire n865;
// (14, 20, 'lutff_3/cout')
// (14, 20, 'lutff_4/in_3')

wire n866;
// (14, 20, 'lutff_4/cout')
// (14, 20, 'lutff_5/in_3')

wire n867;
// (14, 20, 'lutff_5/cout')
// (14, 20, 'lutff_6/in_3')

wire n868;
// (14, 20, 'lutff_6/cout')
// (14, 20, 'lutff_7/in_3')

wire n869;
// (14, 20, 'neigh_op_tnr_0')
// (14, 21, 'neigh_op_rgt_0')
// (14, 22, 'neigh_op_bnr_0')
// (15, 20, 'neigh_op_top_0')
// (15, 21, 'local_g3_0')
// (15, 21, 'lutff_0/in_1')
// (15, 21, 'lutff_0/out')
// (15, 22, 'neigh_op_bot_0')
// (16, 20, 'neigh_op_tnl_0')
// (16, 21, 'neigh_op_lft_0')
// (16, 22, 'neigh_op_bnl_0')

wire n870;
// (14, 20, 'neigh_op_tnr_1')
// (14, 21, 'neigh_op_rgt_1')
// (14, 22, 'neigh_op_bnr_1')
// (15, 20, 'neigh_op_top_1')
// (15, 21, 'local_g3_1')
// (15, 21, 'lutff_1/in_1')
// (15, 21, 'lutff_1/out')
// (15, 22, 'neigh_op_bot_1')
// (16, 20, 'neigh_op_tnl_1')
// (16, 21, 'neigh_op_lft_1')
// (16, 22, 'neigh_op_bnl_1')

wire n871;
// (14, 20, 'neigh_op_tnr_2')
// (14, 21, 'neigh_op_rgt_2')
// (14, 22, 'neigh_op_bnr_2')
// (15, 20, 'neigh_op_top_2')
// (15, 21, 'local_g1_2')
// (15, 21, 'lutff_2/in_1')
// (15, 21, 'lutff_2/out')
// (15, 22, 'neigh_op_bot_2')
// (16, 20, 'neigh_op_tnl_2')
// (16, 21, 'neigh_op_lft_2')
// (16, 22, 'neigh_op_bnl_2')

wire n872;
// (14, 20, 'neigh_op_tnr_3')
// (14, 21, 'neigh_op_rgt_3')
// (14, 22, 'neigh_op_bnr_3')
// (15, 20, 'neigh_op_top_3')
// (15, 21, 'local_g1_3')
// (15, 21, 'lutff_3/in_1')
// (15, 21, 'lutff_3/out')
// (15, 22, 'neigh_op_bot_3')
// (16, 20, 'neigh_op_tnl_3')
// (16, 21, 'neigh_op_lft_3')
// (16, 22, 'neigh_op_bnl_3')

wire n873;
// (14, 20, 'neigh_op_tnr_4')
// (14, 21, 'neigh_op_rgt_4')
// (14, 22, 'neigh_op_bnr_4')
// (15, 20, 'neigh_op_top_4')
// (15, 21, 'local_g3_4')
// (15, 21, 'lutff_4/in_1')
// (15, 21, 'lutff_4/out')
// (15, 22, 'neigh_op_bot_4')
// (16, 20, 'neigh_op_tnl_4')
// (16, 21, 'neigh_op_lft_4')
// (16, 22, 'neigh_op_bnl_4')

wire n874;
// (14, 20, 'neigh_op_tnr_5')
// (14, 21, 'neigh_op_rgt_5')
// (14, 22, 'neigh_op_bnr_5')
// (15, 20, 'neigh_op_top_5')
// (15, 21, 'local_g3_5')
// (15, 21, 'lutff_5/in_1')
// (15, 21, 'lutff_5/out')
// (15, 22, 'neigh_op_bot_5')
// (16, 20, 'neigh_op_tnl_5')
// (16, 21, 'neigh_op_lft_5')
// (16, 22, 'neigh_op_bnl_5')

wire n875;
// (14, 20, 'neigh_op_tnr_6')
// (14, 21, 'neigh_op_rgt_6')
// (14, 22, 'neigh_op_bnr_6')
// (15, 20, 'neigh_op_top_6')
// (15, 21, 'local_g1_6')
// (15, 21, 'lutff_6/in_1')
// (15, 21, 'lutff_6/out')
// (15, 22, 'neigh_op_bot_6')
// (16, 20, 'neigh_op_tnl_6')
// (16, 21, 'neigh_op_lft_6')
// (16, 22, 'neigh_op_bnl_6')

wire n876;
// (14, 20, 'neigh_op_tnr_7')
// (14, 21, 'neigh_op_rgt_7')
// (14, 22, 'neigh_op_bnr_7')
// (15, 20, 'neigh_op_top_7')
// (15, 21, 'local_g1_7')
// (15, 21, 'lutff_7/in_1')
// (15, 21, 'lutff_7/out')
// (15, 22, 'neigh_op_bot_7')
// (16, 20, 'neigh_op_tnl_7')
// (16, 21, 'neigh_op_lft_7')
// (16, 22, 'neigh_op_bnl_7')

reg n877 = 0;
// (14, 20, 'sp4_r_v_b_38')
// (14, 21, 'sp4_r_v_b_27')
// (14, 22, 'sp4_r_v_b_14')
// (14, 23, 'sp4_r_v_b_3')
// (15, 18, 'neigh_op_tnr_2')
// (15, 19, 'neigh_op_rgt_2')
// (15, 19, 'sp4_h_r_9')
// (15, 19, 'sp4_v_t_38')
// (15, 20, 'neigh_op_bnr_2')
// (15, 20, 'sp4_v_b_38')
// (15, 21, 'sp4_v_b_27')
// (15, 22, 'sp4_v_b_14')
// (15, 23, 'sp4_h_r_9')
// (15, 23, 'sp4_v_b_3')
// (16, 18, 'neigh_op_top_2')
// (16, 19, 'lutff_2/out')
// (16, 19, 'sp4_h_r_20')
// (16, 20, 'neigh_op_bot_2')
// (16, 23, 'sp4_h_r_20')
// (17, 18, 'neigh_op_tnl_2')
// (17, 19, 'local_g2_1')
// (17, 19, 'lutff_4/in_1')
// (17, 19, 'neigh_op_lft_2')
// (17, 19, 'sp4_h_r_33')
// (17, 20, 'neigh_op_bnl_2')
// (17, 23, 'local_g2_1')
// (17, 23, 'lutff_4/in_3')
// (17, 23, 'sp4_h_r_33')
// (18, 19, 'sp4_h_r_44')
// (18, 23, 'sp4_h_r_44')
// (19, 19, 'sp4_h_l_44')
// (19, 23, 'sp4_h_l_44')

reg n878 = 0;
// (14, 20, 'sp4_r_v_b_40')
// (14, 21, 'sp4_r_v_b_29')
// (14, 22, 'sp4_r_v_b_16')
// (14, 23, 'sp4_r_v_b_5')
// (15, 18, 'neigh_op_tnr_0')
// (15, 19, 'neigh_op_rgt_0')
// (15, 19, 'sp4_h_r_5')
// (15, 19, 'sp4_v_t_40')
// (15, 20, 'neigh_op_bnr_0')
// (15, 20, 'sp4_v_b_40')
// (15, 21, 'sp4_v_b_29')
// (15, 22, 'sp4_v_b_16')
// (15, 23, 'sp4_h_r_5')
// (15, 23, 'sp4_v_b_5')
// (16, 18, 'neigh_op_top_0')
// (16, 19, 'lutff_0/out')
// (16, 19, 'sp4_h_r_16')
// (16, 20, 'neigh_op_bot_0')
// (16, 23, 'sp4_h_r_16')
// (17, 18, 'neigh_op_tnl_0')
// (17, 19, 'local_g3_5')
// (17, 19, 'lutff_2/in_2')
// (17, 19, 'neigh_op_lft_0')
// (17, 19, 'sp4_h_r_29')
// (17, 20, 'neigh_op_bnl_0')
// (17, 23, 'local_g2_5')
// (17, 23, 'lutff_2/in_3')
// (17, 23, 'sp4_h_r_29')
// (18, 19, 'sp4_h_r_40')
// (18, 23, 'sp4_h_r_40')
// (19, 19, 'sp4_h_l_40')
// (19, 23, 'sp4_h_l_40')

reg io_33_21_1 = 0;
// (14, 21, 'sp12_h_r_0')
// (15, 21, 'sp12_h_r_3')
// (16, 21, 'sp12_h_r_4')
// (17, 20, 'neigh_op_tnr_0')
// (17, 21, 'neigh_op_rgt_0')
// (17, 21, 'sp12_h_r_7')
// (17, 22, 'neigh_op_bnr_0')
// (18, 20, 'neigh_op_top_0')
// (18, 21, 'lutff_0/out')
// (18, 21, 'sp12_h_r_8')
// (18, 22, 'neigh_op_bot_0')
// (19, 20, 'neigh_op_tnl_0')
// (19, 21, 'neigh_op_lft_0')
// (19, 21, 'sp12_h_r_11')
// (19, 22, 'neigh_op_bnl_0')
// (20, 21, 'sp12_h_r_12')
// (21, 21, 'sp12_h_r_15')
// (22, 21, 'sp12_h_r_16')
// (23, 21, 'sp12_h_r_19')
// (24, 21, 'sp12_h_r_20')
// (25, 21, 'sp12_h_r_23')
// (26, 21, 'sp12_h_l_23')
// (26, 21, 'sp12_h_r_0')
// (27, 21, 'sp12_h_r_3')
// (28, 21, 'sp12_h_r_4')
// (29, 21, 'sp12_h_r_7')
// (30, 21, 'sp12_h_r_8')
// (31, 21, 'sp12_h_r_11')
// (32, 21, 'sp12_h_r_12')
// (33, 21, 'io_1/D_OUT_0')
// (33, 21, 'io_1/PAD')
// (33, 21, 'local_g1_4')
// (33, 21, 'span12_horz_12')

wire n880;
// (14, 22, 'sp12_h_r_0')
// (15, 22, 'sp12_h_r_3')
// (16, 22, 'sp12_h_r_4')
// (17, 22, 'sp12_h_r_7')
// (18, 19, 'sp4_r_v_b_37')
// (18, 20, 'sp4_r_v_b_24')
// (18, 21, 'sp4_r_v_b_13')
// (18, 22, 'sp12_h_r_8')
// (18, 22, 'sp4_r_v_b_0')
// (19, 18, 'sp4_v_t_37')
// (19, 19, 'sp4_v_b_37')
// (19, 20, 'sp4_v_b_24')
// (19, 21, 'local_g0_5')
// (19, 21, 'lutff_1/in_2')
// (19, 21, 'sp4_v_b_13')
// (19, 22, 'sp12_h_r_11')
// (19, 22, 'sp4_h_r_7')
// (19, 22, 'sp4_v_b_0')
// (20, 22, 'sp12_h_r_12')
// (20, 22, 'sp4_h_r_18')
// (21, 22, 'sp12_h_r_15')
// (21, 22, 'sp4_h_r_31')
// (22, 22, 'sp12_h_r_16')
// (22, 22, 'sp4_h_r_42')
// (23, 22, 'sp12_h_r_19')
// (23, 22, 'sp4_h_l_42')
// (24, 22, 'sp12_h_r_20')
// (25, 22, 'sp12_h_r_23')
// (26, 10, 'sp12_h_r_0')
// (26, 10, 'sp12_v_t_23')
// (26, 11, 'sp12_v_b_23')
// (26, 12, 'sp12_v_b_20')
// (26, 13, 'sp12_v_b_19')
// (26, 14, 'sp12_v_b_16')
// (26, 15, 'sp12_v_b_15')
// (26, 16, 'sp12_v_b_12')
// (26, 17, 'sp12_v_b_11')
// (26, 18, 'sp12_v_b_8')
// (26, 19, 'sp12_v_b_7')
// (26, 20, 'sp12_v_b_4')
// (26, 21, 'sp12_v_b_3')
// (26, 22, 'sp12_h_l_23')
// (26, 22, 'sp12_v_b_0')
// (27, 10, 'sp12_h_r_3')
// (28, 10, 'sp12_h_r_4')
// (29, 10, 'sp12_h_r_7')
// (30, 10, 'sp12_h_r_8')
// (31, 10, 'sp12_h_r_11')
// (32, 9, 'neigh_op_tnr_2')
// (32, 9, 'neigh_op_tnr_6')
// (32, 10, 'neigh_op_rgt_2')
// (32, 10, 'neigh_op_rgt_6')
// (32, 10, 'sp12_h_r_12')
// (32, 11, 'neigh_op_bnr_2')
// (32, 11, 'neigh_op_bnr_6')
// (33, 10, 'io_1/D_IN_0')
// (33, 10, 'span12_horz_12')

wire n881;
// (14, 22, 'sp4_h_r_3')
// (15, 22, 'sp4_h_r_14')
// (16, 22, 'local_g3_3')
// (16, 22, 'lutff_global/cen')
// (16, 22, 'sp4_h_r_27')
// (17, 19, 'sp4_r_v_b_43')
// (17, 20, 'sp4_r_v_b_30')
// (17, 21, 'neigh_op_tnr_0')
// (17, 21, 'sp4_r_v_b_19')
// (17, 22, 'neigh_op_rgt_0')
// (17, 22, 'sp4_h_r_38')
// (17, 22, 'sp4_r_v_b_6')
// (17, 23, 'neigh_op_bnr_0')
// (17, 23, 'sp4_r_v_b_43')
// (17, 24, 'sp4_r_v_b_30')
// (17, 25, 'sp4_r_v_b_19')
// (17, 26, 'sp4_r_v_b_6')
// (18, 18, 'sp4_v_t_43')
// (18, 19, 'sp4_v_b_43')
// (18, 20, 'sp4_v_b_30')
// (18, 21, 'local_g1_3')
// (18, 21, 'lutff_global/cen')
// (18, 21, 'neigh_op_top_0')
// (18, 21, 'sp4_v_b_19')
// (18, 22, 'lutff_0/out')
// (18, 22, 'sp4_h_l_38')
// (18, 22, 'sp4_h_r_0')
// (18, 22, 'sp4_v_b_6')
// (18, 22, 'sp4_v_t_43')
// (18, 23, 'local_g3_3')
// (18, 23, 'lutff_global/cen')
// (18, 23, 'neigh_op_bot_0')
// (18, 23, 'sp4_v_b_43')
// (18, 24, 'sp4_v_b_30')
// (18, 25, 'sp4_v_b_19')
// (18, 26, 'sp4_v_b_6')
// (19, 21, 'neigh_op_tnl_0')
// (19, 22, 'neigh_op_lft_0')
// (19, 22, 'sp4_h_r_13')
// (19, 23, 'neigh_op_bnl_0')
// (20, 22, 'sp4_h_r_24')
// (21, 22, 'sp4_h_r_37')
// (22, 22, 'sp4_h_l_37')

reg n882 = 0;
// (14, 22, 'sp4_r_v_b_41')
// (14, 23, 'sp4_r_v_b_28')
// (14, 24, 'sp4_r_v_b_17')
// (14, 25, 'neigh_op_tnr_2')
// (14, 25, 'sp4_r_v_b_4')
// (14, 26, 'neigh_op_rgt_2')
// (14, 26, 'sp4_r_v_b_36')
// (14, 27, 'neigh_op_bnr_2')
// (14, 27, 'sp4_r_v_b_25')
// (14, 28, 'sp4_r_v_b_12')
// (14, 29, 'sp4_r_v_b_1')
// (15, 21, 'sp4_h_r_9')
// (15, 21, 'sp4_v_t_41')
// (15, 22, 'sp4_v_b_41')
// (15, 23, 'sp4_v_b_28')
// (15, 24, 'sp4_v_b_17')
// (15, 25, 'neigh_op_top_2')
// (15, 25, 'sp4_v_b_4')
// (15, 25, 'sp4_v_t_36')
// (15, 26, 'local_g3_2')
// (15, 26, 'lutff_2/in_1')
// (15, 26, 'lutff_2/out')
// (15, 26, 'sp4_v_b_36')
// (15, 27, 'neigh_op_bot_2')
// (15, 27, 'sp4_v_b_25')
// (15, 28, 'sp4_v_b_12')
// (15, 29, 'sp4_v_b_1')
// (16, 21, 'sp4_h_r_20')
// (16, 25, 'neigh_op_tnl_2')
// (16, 26, 'neigh_op_lft_2')
// (16, 27, 'neigh_op_bnl_2')
// (17, 21, 'sp4_h_r_33')
// (18, 21, 'local_g3_4')
// (18, 21, 'lutff_2/in_3')
// (18, 21, 'sp4_h_r_44')
// (19, 21, 'sp4_h_l_44')

reg n883 = 0;
// (14, 22, 'sp4_r_v_b_42')
// (14, 23, 'neigh_op_tnr_1')
// (14, 23, 'sp4_r_v_b_31')
// (14, 24, 'neigh_op_rgt_1')
// (14, 24, 'sp4_r_v_b_18')
// (14, 25, 'neigh_op_bnr_1')
// (14, 25, 'sp4_r_v_b_7')
// (15, 21, 'sp4_h_r_0')
// (15, 21, 'sp4_v_t_42')
// (15, 22, 'sp4_v_b_42')
// (15, 23, 'neigh_op_top_1')
// (15, 23, 'sp4_v_b_31')
// (15, 24, 'local_g3_1')
// (15, 24, 'lutff_1/in_1')
// (15, 24, 'lutff_1/out')
// (15, 24, 'sp4_v_b_18')
// (15, 25, 'neigh_op_bot_1')
// (15, 25, 'sp4_v_b_7')
// (16, 21, 'sp4_h_r_13')
// (16, 23, 'neigh_op_tnl_1')
// (16, 24, 'neigh_op_lft_1')
// (16, 25, 'neigh_op_bnl_1')
// (17, 21, 'sp4_h_r_24')
// (18, 21, 'local_g3_5')
// (18, 21, 'lutff_7/in_3')
// (18, 21, 'sp4_h_r_37')
// (19, 21, 'sp4_h_l_37')

reg n884 = 0;
// (14, 22, 'sp4_r_v_b_44')
// (14, 23, 'neigh_op_tnr_2')
// (14, 23, 'sp4_r_v_b_33')
// (14, 24, 'neigh_op_rgt_2')
// (14, 24, 'sp4_r_v_b_20')
// (14, 25, 'neigh_op_bnr_2')
// (14, 25, 'sp4_r_v_b_9')
// (15, 21, 'sp4_h_r_2')
// (15, 21, 'sp4_v_t_44')
// (15, 22, 'sp4_v_b_44')
// (15, 23, 'neigh_op_top_2')
// (15, 23, 'sp4_v_b_33')
// (15, 24, 'local_g1_2')
// (15, 24, 'lutff_2/in_1')
// (15, 24, 'lutff_2/out')
// (15, 24, 'sp4_v_b_20')
// (15, 25, 'neigh_op_bot_2')
// (15, 25, 'sp4_v_b_9')
// (16, 21, 'sp4_h_r_15')
// (16, 23, 'neigh_op_tnl_2')
// (16, 24, 'neigh_op_lft_2')
// (16, 25, 'neigh_op_bnl_2')
// (17, 21, 'sp4_h_r_26')
// (18, 21, 'local_g2_7')
// (18, 21, 'lutff_3/in_0')
// (18, 21, 'sp4_h_r_39')
// (19, 21, 'sp4_h_l_39')

reg n885 = 0;
// (14, 22, 'sp4_r_v_b_47')
// (14, 23, 'sp4_r_v_b_34')
// (14, 24, 'neigh_op_tnr_5')
// (14, 24, 'sp4_r_v_b_23')
// (14, 25, 'neigh_op_rgt_5')
// (14, 25, 'sp4_r_v_b_10')
// (14, 26, 'neigh_op_bnr_5')
// (15, 21, 'sp4_h_r_10')
// (15, 21, 'sp4_v_t_47')
// (15, 22, 'sp4_v_b_47')
// (15, 23, 'sp4_v_b_34')
// (15, 24, 'neigh_op_top_5')
// (15, 24, 'sp4_v_b_23')
// (15, 25, 'local_g1_5')
// (15, 25, 'lutff_5/in_1')
// (15, 25, 'lutff_5/out')
// (15, 25, 'sp4_v_b_10')
// (15, 26, 'neigh_op_bot_5')
// (16, 21, 'sp4_h_r_23')
// (16, 24, 'neigh_op_tnl_5')
// (16, 25, 'neigh_op_lft_5')
// (16, 26, 'neigh_op_bnl_5')
// (17, 21, 'sp4_h_r_34')
// (18, 21, 'local_g3_7')
// (18, 21, 'lutff_4/in_2')
// (18, 21, 'sp4_h_r_47')
// (19, 21, 'sp4_h_l_47')

reg n886 = 0;
// (14, 23, 'neigh_op_tnr_0')
// (14, 24, 'neigh_op_rgt_0')
// (14, 24, 'sp4_h_r_5')
// (14, 25, 'neigh_op_bnr_0')
// (15, 23, 'neigh_op_top_0')
// (15, 24, 'local_g3_0')
// (15, 24, 'lutff_0/in_1')
// (15, 24, 'lutff_0/out')
// (15, 24, 'sp4_h_r_16')
// (15, 25, 'neigh_op_bot_0')
// (16, 23, 'neigh_op_tnl_0')
// (16, 24, 'neigh_op_lft_0')
// (16, 24, 'sp4_h_r_29')
// (16, 25, 'neigh_op_bnl_0')
// (17, 21, 'sp4_r_v_b_40')
// (17, 22, 'sp4_r_v_b_29')
// (17, 23, 'sp4_r_v_b_16')
// (17, 24, 'sp4_h_r_40')
// (17, 24, 'sp4_r_v_b_5')
// (18, 20, 'sp4_v_t_40')
// (18, 21, 'sp4_v_b_40')
// (18, 22, 'sp4_v_b_29')
// (18, 23, 'local_g0_0')
// (18, 23, 'lutff_0/in_2')
// (18, 23, 'sp4_v_b_16')
// (18, 24, 'sp4_h_l_40')
// (18, 24, 'sp4_v_b_5')

reg n887 = 0;
// (14, 23, 'neigh_op_tnr_3')
// (14, 24, 'neigh_op_rgt_3')
// (14, 24, 'sp4_r_v_b_38')
// (14, 25, 'neigh_op_bnr_3')
// (14, 25, 'sp4_r_v_b_27')
// (14, 26, 'sp4_r_v_b_14')
// (14, 27, 'sp4_r_v_b_3')
// (15, 23, 'neigh_op_top_3')
// (15, 23, 'sp4_h_r_3')
// (15, 23, 'sp4_v_t_38')
// (15, 24, 'local_g1_3')
// (15, 24, 'lutff_3/in_1')
// (15, 24, 'lutff_3/out')
// (15, 24, 'sp4_v_b_38')
// (15, 25, 'neigh_op_bot_3')
// (15, 25, 'sp4_v_b_27')
// (15, 26, 'sp4_v_b_14')
// (15, 27, 'sp4_v_b_3')
// (16, 23, 'neigh_op_tnl_3')
// (16, 23, 'sp4_h_r_14')
// (16, 24, 'neigh_op_lft_3')
// (16, 25, 'neigh_op_bnl_3')
// (17, 23, 'sp4_h_r_27')
// (18, 23, 'local_g2_6')
// (18, 23, 'lutff_5/in_1')
// (18, 23, 'sp4_h_r_38')
// (19, 23, 'sp4_h_l_38')

reg n888 = 0;
// (14, 23, 'neigh_op_tnr_4')
// (14, 24, 'neigh_op_rgt_4')
// (14, 25, 'neigh_op_bnr_4')
// (15, 22, 'sp4_r_v_b_46')
// (15, 23, 'neigh_op_top_4')
// (15, 23, 'sp4_r_v_b_35')
// (15, 24, 'local_g3_4')
// (15, 24, 'lutff_4/in_1')
// (15, 24, 'lutff_4/out')
// (15, 24, 'sp4_r_v_b_22')
// (15, 24, 'sp4_r_v_b_41')
// (15, 25, 'neigh_op_bot_4')
// (15, 25, 'sp4_r_v_b_11')
// (15, 25, 'sp4_r_v_b_28')
// (15, 26, 'sp4_r_v_b_17')
// (15, 26, 'sp4_r_v_b_38')
// (15, 27, 'sp4_r_v_b_27')
// (15, 27, 'sp4_r_v_b_4')
// (15, 28, 'sp4_r_v_b_14')
// (15, 28, 'sp4_r_v_b_42')
// (15, 29, 'sp4_r_v_b_3')
// (15, 29, 'sp4_r_v_b_31')
// (15, 30, 'sp4_r_v_b_18')
// (15, 30, 'sp4_r_v_b_42')
// (15, 31, 'sp4_r_v_b_31')
// (15, 31, 'sp4_r_v_b_7')
// (15, 32, 'sp4_r_v_b_18')
// (15, 32, 'sp4_r_v_b_42')
// (16, 21, 'sp4_h_r_4')
// (16, 21, 'sp4_v_t_46')
// (16, 22, 'sp4_v_b_46')
// (16, 23, 'neigh_op_tnl_4')
// (16, 23, 'sp4_v_b_35')
// (16, 23, 'sp4_v_t_41')
// (16, 24, 'neigh_op_lft_4')
// (16, 24, 'sp4_v_b_22')
// (16, 24, 'sp4_v_b_41')
// (16, 25, 'neigh_op_bnl_4')
// (16, 25, 'sp4_v_b_11')
// (16, 25, 'sp4_v_b_28')
// (16, 25, 'sp4_v_t_38')
// (16, 26, 'sp4_v_b_17')
// (16, 26, 'sp4_v_b_38')
// (16, 27, 'sp4_v_b_27')
// (16, 27, 'sp4_v_b_4')
// (16, 27, 'sp4_v_t_42')
// (16, 28, 'sp4_v_b_14')
// (16, 28, 'sp4_v_b_42')
// (16, 29, 'sp4_v_b_3')
// (16, 29, 'sp4_v_b_31')
// (16, 29, 'sp4_v_t_42')
// (16, 30, 'sp4_v_b_18')
// (16, 30, 'sp4_v_b_42')
// (16, 31, 'sp4_v_b_31')
// (16, 31, 'sp4_v_b_7')
// (16, 31, 'sp4_v_t_42')
// (16, 32, 'sp4_v_b_18')
// (16, 32, 'sp4_v_b_42')
// (16, 33, 'span4_vert_31')
// (16, 33, 'span4_vert_7')
// (17, 21, 'sp4_h_r_17')
// (18, 21, 'local_g2_4')
// (18, 21, 'lutff_5/in_3')
// (18, 21, 'sp4_h_r_28')
// (19, 21, 'sp4_h_r_41')
// (20, 21, 'sp4_h_l_41')

reg n889 = 0;
// (14, 23, 'neigh_op_tnr_5')
// (14, 24, 'neigh_op_rgt_5')
// (14, 24, 'sp4_r_v_b_42')
// (14, 25, 'neigh_op_bnr_5')
// (14, 25, 'sp4_r_v_b_31')
// (14, 26, 'sp4_r_v_b_18')
// (14, 27, 'sp4_r_v_b_7')
// (15, 23, 'neigh_op_top_5')
// (15, 23, 'sp4_h_r_0')
// (15, 23, 'sp4_v_t_42')
// (15, 24, 'local_g1_5')
// (15, 24, 'lutff_5/in_1')
// (15, 24, 'lutff_5/out')
// (15, 24, 'sp4_v_b_42')
// (15, 25, 'neigh_op_bot_5')
// (15, 25, 'sp4_v_b_31')
// (15, 26, 'sp4_v_b_18')
// (15, 27, 'sp4_v_b_7')
// (16, 23, 'neigh_op_tnl_5')
// (16, 23, 'sp4_h_r_13')
// (16, 24, 'neigh_op_lft_5')
// (16, 25, 'neigh_op_bnl_5')
// (17, 23, 'sp4_h_r_24')
// (18, 23, 'local_g3_5')
// (18, 23, 'lutff_4/in_0')
// (18, 23, 'sp4_h_r_37')
// (19, 23, 'sp4_h_l_37')

reg n890 = 0;
// (14, 23, 'neigh_op_tnr_6')
// (14, 24, 'neigh_op_rgt_6')
// (14, 24, 'sp4_r_v_b_44')
// (14, 25, 'neigh_op_bnr_6')
// (14, 25, 'sp4_r_v_b_33')
// (14, 26, 'sp4_r_v_b_20')
// (14, 27, 'sp4_r_v_b_9')
// (15, 23, 'neigh_op_top_6')
// (15, 23, 'sp4_h_r_2')
// (15, 23, 'sp4_v_t_44')
// (15, 24, 'local_g1_6')
// (15, 24, 'lutff_6/in_1')
// (15, 24, 'lutff_6/out')
// (15, 24, 'sp4_v_b_44')
// (15, 25, 'neigh_op_bot_6')
// (15, 25, 'sp4_v_b_33')
// (15, 26, 'sp4_v_b_20')
// (15, 27, 'sp4_v_b_9')
// (16, 23, 'neigh_op_tnl_6')
// (16, 23, 'sp4_h_r_15')
// (16, 24, 'neigh_op_lft_6')
// (16, 25, 'neigh_op_bnl_6')
// (17, 23, 'sp4_h_r_26')
// (18, 23, 'local_g2_7')
// (18, 23, 'lutff_1/in_0')
// (18, 23, 'sp4_h_r_39')
// (19, 23, 'sp4_h_l_39')

reg n891 = 0;
// (14, 23, 'neigh_op_tnr_7')
// (14, 24, 'neigh_op_rgt_7')
// (14, 25, 'neigh_op_bnr_7')
// (15, 22, 'sp4_r_v_b_39')
// (15, 23, 'neigh_op_top_7')
// (15, 23, 'sp4_r_v_b_26')
// (15, 24, 'local_g3_7')
// (15, 24, 'lutff_7/in_1')
// (15, 24, 'lutff_7/out')
// (15, 24, 'sp4_r_v_b_15')
// (15, 25, 'neigh_op_bot_7')
// (15, 25, 'sp4_r_v_b_2')
// (16, 21, 'sp4_v_t_39')
// (16, 22, 'local_g3_7')
// (16, 22, 'lutff_0/in_2')
// (16, 22, 'sp4_v_b_39')
// (16, 23, 'neigh_op_tnl_7')
// (16, 23, 'sp4_v_b_26')
// (16, 24, 'neigh_op_lft_7')
// (16, 24, 'sp4_v_b_15')
// (16, 25, 'neigh_op_bnl_7')
// (16, 25, 'sp4_v_b_2')

reg n892 = 0;
// (14, 23, 'sp4_r_v_b_42')
// (14, 24, 'neigh_op_tnr_1')
// (14, 24, 'sp4_r_v_b_31')
// (14, 25, 'neigh_op_rgt_1')
// (14, 25, 'sp4_r_v_b_18')
// (14, 26, 'neigh_op_bnr_1')
// (14, 26, 'sp4_r_v_b_7')
// (15, 22, 'sp4_h_r_0')
// (15, 22, 'sp4_v_t_42')
// (15, 23, 'sp4_v_b_42')
// (15, 24, 'neigh_op_top_1')
// (15, 24, 'sp4_v_b_31')
// (15, 25, 'local_g3_1')
// (15, 25, 'lutff_1/in_1')
// (15, 25, 'lutff_1/out')
// (15, 25, 'sp4_v_b_18')
// (15, 26, 'neigh_op_bot_1')
// (15, 26, 'sp4_v_b_7')
// (16, 22, 'local_g1_5')
// (16, 22, 'lutff_2/in_2')
// (16, 22, 'sp4_h_r_13')
// (16, 24, 'neigh_op_tnl_1')
// (16, 25, 'neigh_op_lft_1')
// (16, 26, 'neigh_op_bnl_1')
// (17, 22, 'sp4_h_r_24')
// (18, 22, 'sp4_h_r_37')
// (19, 22, 'sp4_h_l_37')

reg n893 = 0;
// (14, 24, 'neigh_op_tnr_0')
// (14, 25, 'neigh_op_rgt_0')
// (14, 26, 'neigh_op_bnr_0')
// (15, 23, 'sp4_r_v_b_41')
// (15, 24, 'neigh_op_top_0')
// (15, 24, 'sp4_r_v_b_28')
// (15, 25, 'local_g3_0')
// (15, 25, 'lutff_0/in_1')
// (15, 25, 'lutff_0/out')
// (15, 25, 'sp4_r_v_b_17')
// (15, 26, 'neigh_op_bot_0')
// (15, 26, 'sp4_r_v_b_4')
// (16, 22, 'local_g1_4')
// (16, 22, 'lutff_1/in_0')
// (16, 22, 'sp4_h_r_4')
// (16, 22, 'sp4_v_t_41')
// (16, 23, 'sp4_v_b_41')
// (16, 24, 'neigh_op_tnl_0')
// (16, 24, 'sp4_v_b_28')
// (16, 25, 'neigh_op_lft_0')
// (16, 25, 'sp4_v_b_17')
// (16, 26, 'neigh_op_bnl_0')
// (16, 26, 'sp4_v_b_4')
// (17, 22, 'sp4_h_r_17')
// (18, 22, 'sp4_h_r_28')
// (19, 22, 'sp4_h_r_41')
// (20, 22, 'sp4_h_l_41')

reg n894 = 0;
// (14, 24, 'neigh_op_tnr_2')
// (14, 25, 'neigh_op_rgt_2')
// (14, 25, 'sp4_h_r_9')
// (14, 26, 'neigh_op_bnr_2')
// (15, 24, 'neigh_op_top_2')
// (15, 25, 'local_g1_2')
// (15, 25, 'lutff_2/in_1')
// (15, 25, 'lutff_2/out')
// (15, 25, 'sp4_h_r_20')
// (15, 26, 'neigh_op_bot_2')
// (16, 24, 'neigh_op_tnl_2')
// (16, 25, 'neigh_op_lft_2')
// (16, 25, 'sp4_h_r_33')
// (16, 26, 'neigh_op_bnl_2')
// (17, 22, 'sp4_r_v_b_44')
// (17, 23, 'sp4_r_v_b_33')
// (17, 24, 'sp4_r_v_b_20')
// (17, 25, 'sp4_h_r_44')
// (17, 25, 'sp4_r_v_b_9')
// (18, 21, 'sp4_v_t_44')
// (18, 22, 'sp4_v_b_44')
// (18, 23, 'local_g2_1')
// (18, 23, 'lutff_2/in_1')
// (18, 23, 'sp4_v_b_33')
// (18, 24, 'sp4_v_b_20')
// (18, 25, 'sp4_h_l_44')
// (18, 25, 'sp4_v_b_9')

reg n895 = 0;
// (14, 24, 'neigh_op_tnr_3')
// (14, 25, 'neigh_op_rgt_3')
// (14, 25, 'sp4_h_r_11')
// (14, 26, 'neigh_op_bnr_3')
// (15, 24, 'neigh_op_top_3')
// (15, 25, 'local_g1_3')
// (15, 25, 'lutff_3/in_1')
// (15, 25, 'lutff_3/out')
// (15, 25, 'sp4_h_r_22')
// (15, 26, 'neigh_op_bot_3')
// (16, 24, 'neigh_op_tnl_3')
// (16, 25, 'neigh_op_lft_3')
// (16, 25, 'sp4_h_r_35')
// (16, 26, 'neigh_op_bnl_3')
// (17, 22, 'sp4_r_v_b_37')
// (17, 23, 'sp4_r_v_b_24')
// (17, 24, 'sp4_r_v_b_13')
// (17, 25, 'sp4_h_r_46')
// (17, 25, 'sp4_r_v_b_0')
// (17, 26, 'sp4_r_v_b_41')
// (17, 27, 'sp4_r_v_b_28')
// (17, 28, 'sp4_r_v_b_17')
// (17, 29, 'sp4_r_v_b_4')
// (18, 21, 'sp4_v_t_37')
// (18, 22, 'sp4_v_b_37')
// (18, 23, 'local_g2_0')
// (18, 23, 'lutff_3/in_3')
// (18, 23, 'sp4_v_b_24')
// (18, 24, 'sp4_v_b_13')
// (18, 25, 'sp4_h_l_46')
// (18, 25, 'sp4_v_b_0')
// (18, 25, 'sp4_v_t_41')
// (18, 26, 'sp4_v_b_41')
// (18, 27, 'sp4_v_b_28')
// (18, 28, 'sp4_v_b_17')
// (18, 29, 'sp4_v_b_4')

reg n896 = 0;
// (14, 24, 'neigh_op_tnr_6')
// (14, 24, 'sp4_r_v_b_41')
// (14, 25, 'neigh_op_rgt_6')
// (14, 25, 'sp4_r_v_b_28')
// (14, 26, 'neigh_op_bnr_6')
// (14, 26, 'sp4_r_v_b_17')
// (14, 27, 'sp4_r_v_b_4')
// (15, 23, 'sp4_h_r_4')
// (15, 23, 'sp4_v_t_41')
// (15, 24, 'neigh_op_top_6')
// (15, 24, 'sp4_v_b_41')
// (15, 25, 'local_g1_6')
// (15, 25, 'lutff_6/in_1')
// (15, 25, 'lutff_6/out')
// (15, 25, 'sp4_v_b_28')
// (15, 26, 'neigh_op_bot_6')
// (15, 26, 'sp4_v_b_17')
// (15, 27, 'sp4_v_b_4')
// (16, 23, 'sp4_h_r_17')
// (16, 24, 'neigh_op_tnl_6')
// (16, 25, 'neigh_op_lft_6')
// (16, 26, 'neigh_op_bnl_6')
// (17, 23, 'sp4_h_r_28')
// (18, 23, 'local_g3_1')
// (18, 23, 'lutff_6/in_2')
// (18, 23, 'sp4_h_r_41')
// (19, 23, 'sp4_h_l_41')

reg n897 = 0;
// (14, 24, 'neigh_op_tnr_7')
// (14, 25, 'neigh_op_rgt_7')
// (14, 26, 'neigh_op_bnr_7')
// (15, 24, 'neigh_op_top_7')
// (15, 24, 'sp4_r_v_b_42')
// (15, 25, 'local_g1_7')
// (15, 25, 'lutff_7/in_1')
// (15, 25, 'lutff_7/out')
// (15, 25, 'sp4_r_v_b_31')
// (15, 26, 'neigh_op_bot_7')
// (15, 26, 'sp4_r_v_b_18')
// (15, 27, 'sp4_r_v_b_7')
// (16, 23, 'sp4_h_r_7')
// (16, 23, 'sp4_v_t_42')
// (16, 24, 'neigh_op_tnl_7')
// (16, 24, 'sp4_v_b_42')
// (16, 25, 'neigh_op_lft_7')
// (16, 25, 'sp4_v_b_31')
// (16, 26, 'neigh_op_bnl_7')
// (16, 26, 'sp4_v_b_18')
// (16, 27, 'sp4_v_b_7')
// (17, 23, 'sp4_h_r_18')
// (18, 23, 'local_g3_7')
// (18, 23, 'lutff_7/in_3')
// (18, 23, 'sp4_h_r_31')
// (19, 23, 'sp4_h_r_42')
// (20, 23, 'sp4_h_l_42')

reg n898 = 0;
// (14, 24, 'sp4_r_v_b_40')
// (14, 25, 'neigh_op_tnr_0')
// (14, 25, 'sp4_r_v_b_29')
// (14, 26, 'neigh_op_rgt_0')
// (14, 26, 'sp4_r_v_b_16')
// (14, 27, 'neigh_op_bnr_0')
// (14, 27, 'sp4_r_v_b_5')
// (15, 23, 'sp4_h_r_10')
// (15, 23, 'sp4_v_t_40')
// (15, 24, 'sp4_v_b_40')
// (15, 25, 'neigh_op_top_0')
// (15, 25, 'sp4_v_b_29')
// (15, 26, 'local_g3_0')
// (15, 26, 'lutff_0/in_1')
// (15, 26, 'lutff_0/out')
// (15, 26, 'sp4_v_b_16')
// (15, 27, 'neigh_op_bot_0')
// (15, 27, 'sp4_v_b_5')
// (16, 23, 'sp4_h_r_23')
// (16, 25, 'neigh_op_tnl_0')
// (16, 26, 'neigh_op_lft_0')
// (16, 27, 'neigh_op_bnl_0')
// (17, 23, 'sp4_h_r_34')
// (18, 20, 'sp4_r_v_b_47')
// (18, 21, 'local_g2_2')
// (18, 21, 'lutff_0/in_0')
// (18, 21, 'sp4_r_v_b_34')
// (18, 22, 'sp4_r_v_b_23')
// (18, 23, 'sp4_h_r_47')
// (18, 23, 'sp4_r_v_b_10')
// (19, 19, 'sp4_v_t_47')
// (19, 20, 'sp4_v_b_47')
// (19, 21, 'sp4_v_b_34')
// (19, 22, 'sp4_v_b_23')
// (19, 23, 'sp4_h_l_47')
// (19, 23, 'sp4_v_b_10')

reg n899 = 0;
// (14, 25, 'neigh_op_tnr_1')
// (14, 25, 'sp4_r_v_b_47')
// (14, 26, 'neigh_op_rgt_1')
// (14, 26, 'sp4_r_v_b_34')
// (14, 27, 'neigh_op_bnr_1')
// (14, 27, 'sp4_r_v_b_23')
// (14, 28, 'sp4_r_v_b_10')
// (15, 24, 'sp4_h_r_10')
// (15, 24, 'sp4_v_t_47')
// (15, 25, 'neigh_op_top_1')
// (15, 25, 'sp4_v_b_47')
// (15, 26, 'local_g3_1')
// (15, 26, 'lutff_1/in_1')
// (15, 26, 'lutff_1/out')
// (15, 26, 'sp4_v_b_34')
// (15, 27, 'neigh_op_bot_1')
// (15, 27, 'sp4_v_b_23')
// (15, 28, 'sp4_v_b_10')
// (16, 24, 'sp4_h_r_23')
// (16, 25, 'neigh_op_tnl_1')
// (16, 26, 'neigh_op_lft_1')
// (16, 27, 'neigh_op_bnl_1')
// (17, 24, 'sp4_h_r_34')
// (18, 21, 'local_g3_3')
// (18, 21, 'lutff_1/in_1')
// (18, 21, 'sp4_r_v_b_43')
// (18, 22, 'sp4_r_v_b_30')
// (18, 23, 'sp4_r_v_b_19')
// (18, 24, 'sp4_h_r_47')
// (18, 24, 'sp4_r_v_b_6')
// (19, 20, 'sp4_v_t_43')
// (19, 21, 'sp4_v_b_43')
// (19, 22, 'sp4_v_b_30')
// (19, 23, 'sp4_v_b_19')
// (19, 24, 'sp4_h_l_47')
// (19, 24, 'sp4_h_r_1')
// (19, 24, 'sp4_v_b_6')
// (20, 24, 'sp4_h_r_12')
// (21, 24, 'sp4_h_r_25')
// (22, 24, 'sp4_h_r_36')
// (23, 24, 'sp4_h_l_36')

reg n900 = 0;
// (15, 6, 'neigh_op_tnr_0')
// (15, 7, 'local_g3_0')
// (15, 7, 'lutff_3/in_2')
// (15, 7, 'neigh_op_rgt_0')
// (15, 8, 'neigh_op_bnr_0')
// (16, 6, 'neigh_op_top_0')
// (16, 7, 'local_g3_0')
// (16, 7, 'lutff_0/in_1')
// (16, 7, 'lutff_0/out')
// (16, 8, 'neigh_op_bot_0')
// (17, 6, 'neigh_op_tnl_0')
// (17, 7, 'neigh_op_lft_0')
// (17, 8, 'neigh_op_bnl_0')

reg n901 = 0;
// (15, 6, 'neigh_op_tnr_1')
// (15, 7, 'local_g3_1')
// (15, 7, 'lutff_3/in_1')
// (15, 7, 'neigh_op_rgt_1')
// (15, 8, 'neigh_op_bnr_1')
// (16, 6, 'neigh_op_top_1')
// (16, 7, 'local_g3_1')
// (16, 7, 'lutff_1/in_1')
// (16, 7, 'lutff_1/out')
// (16, 8, 'neigh_op_bot_1')
// (17, 6, 'neigh_op_tnl_1')
// (17, 7, 'neigh_op_lft_1')
// (17, 8, 'neigh_op_bnl_1')

reg n902 = 0;
// (15, 6, 'neigh_op_tnr_2')
// (15, 7, 'local_g2_2')
// (15, 7, 'lutff_0/in_2')
// (15, 7, 'lutff_4/in_0')
// (15, 7, 'neigh_op_rgt_2')
// (15, 8, 'neigh_op_bnr_2')
// (16, 6, 'neigh_op_top_2')
// (16, 7, 'local_g1_2')
// (16, 7, 'lutff_2/in_1')
// (16, 7, 'lutff_2/out')
// (16, 8, 'neigh_op_bot_2')
// (17, 6, 'neigh_op_tnl_2')
// (17, 7, 'neigh_op_lft_2')
// (17, 8, 'neigh_op_bnl_2')

reg n903 = 0;
// (15, 6, 'neigh_op_tnr_3')
// (15, 7, 'local_g2_3')
// (15, 7, 'lutff_3/in_0')
// (15, 7, 'neigh_op_rgt_3')
// (15, 8, 'neigh_op_bnr_3')
// (16, 6, 'neigh_op_top_3')
// (16, 7, 'local_g1_3')
// (16, 7, 'lutff_3/in_1')
// (16, 7, 'lutff_3/out')
// (16, 8, 'neigh_op_bot_3')
// (17, 6, 'neigh_op_tnl_3')
// (17, 7, 'neigh_op_lft_3')
// (17, 8, 'neigh_op_bnl_3')

reg n904 = 0;
// (15, 6, 'neigh_op_tnr_4')
// (15, 7, 'local_g2_4')
// (15, 7, 'lutff_3/in_3')
// (15, 7, 'neigh_op_rgt_4')
// (15, 8, 'neigh_op_bnr_4')
// (16, 6, 'neigh_op_top_4')
// (16, 7, 'local_g3_4')
// (16, 7, 'lutff_4/in_1')
// (16, 7, 'lutff_4/out')
// (16, 8, 'neigh_op_bot_4')
// (17, 6, 'neigh_op_tnl_4')
// (17, 7, 'neigh_op_lft_4')
// (17, 8, 'neigh_op_bnl_4')

reg n905 = 0;
// (15, 6, 'neigh_op_tnr_5')
// (15, 7, 'local_g2_5')
// (15, 7, 'lutff_0/in_1')
// (15, 7, 'lutff_4/in_3')
// (15, 7, 'neigh_op_rgt_5')
// (15, 8, 'neigh_op_bnr_5')
// (16, 6, 'neigh_op_top_5')
// (16, 7, 'local_g3_5')
// (16, 7, 'lutff_5/in_1')
// (16, 7, 'lutff_5/out')
// (16, 8, 'neigh_op_bot_5')
// (17, 6, 'neigh_op_tnl_5')
// (17, 7, 'neigh_op_lft_5')
// (17, 8, 'neigh_op_bnl_5')

wire n906;
// (15, 7, 'lutff_1/lout')
// (15, 7, 'lutff_2/in_2')

wire n907;
// (15, 7, 'lutff_3/lout')
// (15, 7, 'lutff_4/in_2')

wire n908;
// (15, 7, 'lutff_5/lout')
// (15, 7, 'lutff_6/in_2')

reg n909 = 0;
// (15, 7, 'neigh_op_tnr_6')
// (15, 8, 'neigh_op_rgt_6')
// (15, 8, 'sp4_r_v_b_44')
// (15, 9, 'neigh_op_bnr_6')
// (15, 9, 'sp4_r_v_b_33')
// (15, 10, 'sp4_r_v_b_20')
// (15, 11, 'sp4_r_v_b_9')
// (16, 7, 'neigh_op_top_6')
// (16, 7, 'sp4_v_t_44')
// (16, 8, 'lutff_6/out')
// (16, 8, 'sp4_v_b_44')
// (16, 9, 'neigh_op_bot_6')
// (16, 9, 'sp4_v_b_33')
// (16, 10, 'local_g0_4')
// (16, 10, 'lutff_7/in_3')
// (16, 10, 'sp4_v_b_20')
// (16, 11, 'sp4_v_b_9')
// (17, 7, 'neigh_op_tnl_6')
// (17, 8, 'neigh_op_lft_6')
// (17, 9, 'neigh_op_bnl_6')

reg n910 = 0;
// (15, 8, 'local_g0_2')
// (15, 8, 'lutff_7/in_1')
// (15, 8, 'sp4_h_r_10')
// (16, 7, 'neigh_op_tnr_1')
// (16, 8, 'neigh_op_rgt_1')
// (16, 8, 'sp4_h_r_23')
// (16, 9, 'neigh_op_bnr_1')
// (17, 7, 'neigh_op_top_1')
// (17, 8, 'lutff_1/out')
// (17, 8, 'sp4_h_r_34')
// (17, 9, 'neigh_op_bot_1')
// (18, 7, 'neigh_op_tnl_1')
// (18, 8, 'neigh_op_lft_1')
// (18, 8, 'sp4_h_r_47')
// (18, 9, 'neigh_op_bnl_1')
// (19, 8, 'sp4_h_l_47')

reg n911 = 0;
// (15, 8, 'local_g1_0')
// (15, 8, 'lutff_0/in_1')
// (15, 8, 'sp4_h_r_0')
// (16, 7, 'neigh_op_tnr_4')
// (16, 8, 'neigh_op_rgt_4')
// (16, 8, 'sp4_h_r_13')
// (16, 9, 'neigh_op_bnr_4')
// (17, 7, 'neigh_op_top_4')
// (17, 8, 'lutff_4/out')
// (17, 8, 'sp4_h_r_24')
// (17, 9, 'neigh_op_bot_4')
// (18, 7, 'neigh_op_tnl_4')
// (18, 8, 'neigh_op_lft_4')
// (18, 8, 'sp4_h_r_37')
// (18, 9, 'neigh_op_bnl_4')
// (19, 8, 'sp4_h_l_37')

wire n912;
// (15, 8, 'lutff_0/lout')
// (15, 8, 'lutff_1/in_2')

reg n913 = 0;
// (15, 8, 'neigh_op_tnr_0')
// (15, 9, 'neigh_op_rgt_0')
// (15, 10, 'neigh_op_bnr_0')
// (16, 5, 'sp12_v_t_23')
// (16, 6, 'sp12_v_b_23')
// (16, 7, 'sp12_v_b_20')
// (16, 8, 'neigh_op_top_0')
// (16, 8, 'sp12_v_b_19')
// (16, 9, 'lutff_0/out')
// (16, 9, 'sp12_v_b_16')
// (16, 10, 'neigh_op_bot_0')
// (16, 10, 'sp12_v_b_15')
// (16, 11, 'sp12_v_b_12')
// (16, 12, 'sp12_v_b_11')
// (16, 13, 'sp12_v_b_8')
// (16, 14, 'sp12_v_b_7')
// (16, 15, 'sp12_v_b_4')
// (16, 16, 'sp12_v_b_3')
// (16, 17, 'sp12_h_r_0')
// (16, 17, 'sp12_v_b_0')
// (17, 8, 'neigh_op_tnl_0')
// (17, 9, 'neigh_op_lft_0')
// (17, 10, 'neigh_op_bnl_0')
// (17, 17, 'local_g1_3')
// (17, 17, 'lutff_1/in_3')
// (17, 17, 'sp12_h_r_3')
// (18, 17, 'sp12_h_r_4')
// (19, 17, 'sp12_h_r_7')
// (20, 17, 'sp12_h_r_8')
// (21, 17, 'sp12_h_r_11')
// (22, 17, 'sp12_h_r_12')
// (23, 17, 'sp12_h_r_15')
// (24, 17, 'sp12_h_r_16')
// (25, 17, 'sp12_h_r_19')
// (26, 17, 'sp12_h_r_20')
// (27, 17, 'sp12_h_r_23')
// (28, 17, 'sp12_h_l_23')

reg n914 = 0;
// (15, 8, 'sp4_r_v_b_46')
// (15, 9, 'sp4_r_v_b_35')
// (15, 10, 'sp4_r_v_b_22')
// (15, 11, 'sp4_r_v_b_11')
// (16, 6, 'neigh_op_tnr_0')
// (16, 7, 'neigh_op_rgt_0')
// (16, 7, 'sp4_h_r_5')
// (16, 7, 'sp4_v_t_46')
// (16, 8, 'neigh_op_bnr_0')
// (16, 8, 'sp4_v_b_46')
// (16, 9, 'sp4_v_b_35')
// (16, 10, 'local_g1_6')
// (16, 10, 'lutff_0/in_3')
// (16, 10, 'sp4_v_b_22')
// (16, 11, 'sp4_v_b_11')
// (17, 6, 'neigh_op_top_0')
// (17, 7, 'lutff_0/out')
// (17, 7, 'sp4_h_r_16')
// (17, 8, 'neigh_op_bot_0')
// (18, 6, 'neigh_op_tnl_0')
// (18, 7, 'neigh_op_lft_0')
// (18, 7, 'sp4_h_r_29')
// (18, 8, 'neigh_op_bnl_0')
// (19, 7, 'sp4_h_r_40')
// (20, 7, 'sp4_h_l_40')

reg n915 = 0;
// (15, 9, 'local_g0_1')
// (15, 9, 'lutff_2/in_1')
// (15, 9, 'sp4_h_r_1')
// (16, 9, 'sp4_h_r_12')
// (17, 8, 'neigh_op_tnr_2')
// (17, 9, 'neigh_op_rgt_2')
// (17, 9, 'sp4_h_r_25')
// (17, 10, 'neigh_op_bnr_2')
// (18, 8, 'neigh_op_top_2')
// (18, 9, 'lutff_2/out')
// (18, 9, 'sp4_h_r_36')
// (18, 10, 'neigh_op_bot_2')
// (19, 8, 'neigh_op_tnl_2')
// (19, 9, 'neigh_op_lft_2')
// (19, 9, 'sp4_h_l_36')
// (19, 10, 'neigh_op_bnl_2')

reg n916 = 0;
// (15, 9, 'local_g0_3')
// (15, 9, 'lutff_0/in_3')
// (15, 9, 'sp4_h_r_11')
// (16, 9, 'sp4_h_r_22')
// (17, 8, 'neigh_op_tnr_7')
// (17, 9, 'neigh_op_rgt_7')
// (17, 9, 'sp4_h_r_35')
// (17, 10, 'neigh_op_bnr_7')
// (18, 8, 'neigh_op_top_7')
// (18, 9, 'lutff_7/out')
// (18, 9, 'sp4_h_r_46')
// (18, 10, 'neigh_op_bot_7')
// (19, 8, 'neigh_op_tnl_7')
// (19, 9, 'neigh_op_lft_7')
// (19, 9, 'sp4_h_l_46')
// (19, 10, 'neigh_op_bnl_7')

reg n917 = 0;
// (15, 9, 'local_g1_5')
// (15, 9, 'lutff_1/in_3')
// (15, 9, 'sp4_h_r_5')
// (16, 9, 'sp4_h_r_16')
// (17, 8, 'neigh_op_tnr_4')
// (17, 9, 'neigh_op_rgt_4')
// (17, 9, 'sp4_h_r_29')
// (17, 10, 'neigh_op_bnr_4')
// (18, 8, 'neigh_op_top_4')
// (18, 9, 'lutff_4/out')
// (18, 9, 'sp4_h_r_40')
// (18, 10, 'neigh_op_bot_4')
// (19, 8, 'neigh_op_tnl_4')
// (19, 9, 'neigh_op_lft_4')
// (19, 9, 'sp4_h_l_40')
// (19, 10, 'neigh_op_bnl_4')

reg n918 = 0;
// (15, 9, 'neigh_op_tnr_0')
// (15, 10, 'local_g3_0')
// (15, 10, 'lutff_4/in_3')
// (15, 10, 'neigh_op_rgt_0')
// (15, 11, 'neigh_op_bnr_0')
// (16, 9, 'neigh_op_top_0')
// (16, 10, 'lutff_0/out')
// (16, 11, 'neigh_op_bot_0')
// (17, 9, 'neigh_op_tnl_0')
// (17, 10, 'neigh_op_lft_0')
// (17, 11, 'neigh_op_bnl_0')

reg n919 = 0;
// (15, 9, 'neigh_op_tnr_2')
// (15, 10, 'local_g2_2')
// (15, 10, 'lutff_7/in_3')
// (15, 10, 'neigh_op_rgt_2')
// (15, 11, 'neigh_op_bnr_2')
// (16, 9, 'neigh_op_top_2')
// (16, 10, 'lutff_2/out')
// (16, 11, 'neigh_op_bot_2')
// (17, 9, 'neigh_op_tnl_2')
// (17, 10, 'neigh_op_lft_2')
// (17, 11, 'neigh_op_bnl_2')

reg n920 = 0;
// (15, 9, 'neigh_op_tnr_3')
// (15, 10, 'neigh_op_rgt_3')
// (15, 11, 'local_g1_3')
// (15, 11, 'lutff_5/in_3')
// (15, 11, 'neigh_op_bnr_3')
// (16, 9, 'neigh_op_top_3')
// (16, 10, 'lutff_3/out')
// (16, 11, 'neigh_op_bot_3')
// (17, 9, 'neigh_op_tnl_3')
// (17, 10, 'neigh_op_lft_3')
// (17, 11, 'neigh_op_bnl_3')

reg n921 = 0;
// (15, 9, 'neigh_op_tnr_4')
// (15, 10, 'neigh_op_rgt_4')
// (15, 11, 'local_g1_4')
// (15, 11, 'lutff_6/in_3')
// (15, 11, 'neigh_op_bnr_4')
// (16, 9, 'neigh_op_top_4')
// (16, 10, 'lutff_4/out')
// (16, 11, 'neigh_op_bot_4')
// (17, 9, 'neigh_op_tnl_4')
// (17, 10, 'neigh_op_lft_4')
// (17, 11, 'neigh_op_bnl_4')

reg n922 = 0;
// (15, 9, 'neigh_op_tnr_6')
// (15, 10, 'local_g3_6')
// (15, 10, 'lutff_1/in_0')
// (15, 10, 'neigh_op_rgt_6')
// (15, 11, 'neigh_op_bnr_6')
// (16, 9, 'neigh_op_top_6')
// (16, 10, 'lutff_6/out')
// (16, 11, 'neigh_op_bot_6')
// (17, 9, 'neigh_op_tnl_6')
// (17, 10, 'neigh_op_lft_6')
// (17, 11, 'neigh_op_bnl_6')

reg n923 = 0;
// (15, 10, 'neigh_op_tnr_0')
// (15, 11, 'neigh_op_rgt_0')
// (15, 12, 'neigh_op_bnr_0')
// (16, 10, 'neigh_op_top_0')
// (16, 10, 'sp4_r_v_b_44')
// (16, 11, 'lutff_0/out')
// (16, 11, 'sp4_r_v_b_33')
// (16, 12, 'neigh_op_bot_0')
// (16, 12, 'sp4_r_v_b_20')
// (16, 13, 'sp4_r_v_b_9')
// (16, 14, 'sp4_r_v_b_37')
// (16, 15, 'sp4_r_v_b_24')
// (16, 16, 'sp4_r_v_b_13')
// (16, 17, 'sp4_r_v_b_0')
// (17, 9, 'sp4_v_t_44')
// (17, 10, 'neigh_op_tnl_0')
// (17, 10, 'sp4_v_b_44')
// (17, 11, 'neigh_op_lft_0')
// (17, 11, 'sp4_v_b_33')
// (17, 12, 'neigh_op_bnl_0')
// (17, 12, 'sp4_v_b_20')
// (17, 13, 'sp4_v_b_9')
// (17, 13, 'sp4_v_t_37')
// (17, 14, 'sp4_v_b_37')
// (17, 15, 'sp4_v_b_24')
// (17, 16, 'sp4_v_b_13')
// (17, 17, 'local_g0_0')
// (17, 17, 'lutff_3/in_1')
// (17, 17, 'sp4_v_b_0')

reg n924 = 0;
// (15, 10, 'neigh_op_tnr_1')
// (15, 11, 'neigh_op_rgt_1')
// (15, 12, 'neigh_op_bnr_1')
// (16, 10, 'neigh_op_top_1')
// (16, 10, 'sp4_r_v_b_46')
// (16, 11, 'lutff_1/out')
// (16, 11, 'sp4_r_v_b_35')
// (16, 12, 'neigh_op_bot_1')
// (16, 12, 'sp4_r_v_b_22')
// (16, 13, 'sp4_r_v_b_11')
// (17, 9, 'sp4_v_t_46')
// (17, 10, 'neigh_op_tnl_1')
// (17, 10, 'sp4_v_b_46')
// (17, 11, 'neigh_op_lft_1')
// (17, 11, 'sp4_v_b_35')
// (17, 12, 'neigh_op_bnl_1')
// (17, 12, 'sp4_v_b_22')
// (17, 13, 'sp4_h_r_5')
// (17, 13, 'sp4_v_b_11')
// (18, 13, 'sp4_h_r_16')
// (19, 13, 'sp4_h_r_29')
// (20, 13, 'local_g3_0')
// (20, 13, 'lutff_0/in_1')
// (20, 13, 'sp4_h_r_40')
// (21, 13, 'sp4_h_l_40')

reg n925 = 0;
// (15, 10, 'neigh_op_tnr_2')
// (15, 11, 'neigh_op_rgt_2')
// (15, 12, 'neigh_op_bnr_2')
// (16, 10, 'neigh_op_top_2')
// (16, 11, 'lutff_2/out')
// (16, 11, 'sp4_h_r_4')
// (16, 12, 'neigh_op_bot_2')
// (17, 10, 'neigh_op_tnl_2')
// (17, 11, 'neigh_op_lft_2')
// (17, 11, 'sp4_h_r_17')
// (17, 12, 'neigh_op_bnl_2')
// (18, 11, 'sp4_h_r_28')
// (19, 11, 'sp4_h_r_41')
// (19, 12, 'sp4_r_v_b_41')
// (19, 13, 'sp4_r_v_b_28')
// (19, 14, 'sp4_r_v_b_17')
// (19, 15, 'sp4_r_v_b_4')
// (20, 11, 'sp4_h_l_41')
// (20, 11, 'sp4_v_t_41')
// (20, 12, 'sp4_v_b_41')
// (20, 13, 'local_g3_4')
// (20, 13, 'lutff_6/in_1')
// (20, 13, 'sp4_v_b_28')
// (20, 14, 'sp4_v_b_17')
// (20, 15, 'sp4_v_b_4')

reg n926 = 0;
// (15, 10, 'neigh_op_tnr_5')
// (15, 11, 'neigh_op_rgt_5')
// (15, 12, 'neigh_op_bnr_5')
// (16, 10, 'neigh_op_top_5')
// (16, 11, 'lutff_5/out')
// (16, 12, 'neigh_op_bot_5')
// (17, 10, 'neigh_op_tnl_5')
// (17, 11, 'local_g0_5')
// (17, 11, 'lutff_0/in_1')
// (17, 11, 'neigh_op_lft_5')
// (17, 12, 'neigh_op_bnl_5')

reg n927 = 0;
// (15, 10, 'neigh_op_tnr_6')
// (15, 11, 'neigh_op_rgt_6')
// (15, 12, 'neigh_op_bnr_6')
// (16, 10, 'neigh_op_top_6')
// (16, 11, 'lutff_6/out')
// (16, 12, 'neigh_op_bot_6')
// (17, 10, 'neigh_op_tnl_6')
// (17, 11, 'local_g0_6')
// (17, 11, 'lutff_5/in_1')
// (17, 11, 'neigh_op_lft_6')
// (17, 12, 'neigh_op_bnl_6')

reg n928 = 0;
// (15, 10, 'neigh_op_tnr_7')
// (15, 11, 'neigh_op_rgt_7')
// (15, 12, 'neigh_op_bnr_7')
// (16, 10, 'neigh_op_top_7')
// (16, 11, 'lutff_7/out')
// (16, 12, 'neigh_op_bot_7')
// (17, 10, 'neigh_op_tnl_7')
// (17, 11, 'neigh_op_lft_7')
// (17, 12, 'local_g2_7')
// (17, 12, 'lutff_4/in_1')
// (17, 12, 'neigh_op_bnl_7')

reg n929 = 0;
// (15, 10, 'sp4_h_r_0')
// (16, 10, 'local_g0_5')
// (16, 10, 'lutff_6/in_3')
// (16, 10, 'sp4_h_r_13')
// (17, 10, 'sp4_h_r_24')
// (18, 10, 'sp4_h_r_37')
// (18, 11, 'sp4_r_v_b_37')
// (18, 12, 'sp4_r_v_b_24')
// (18, 13, 'sp4_r_v_b_13')
// (18, 14, 'sp4_r_v_b_0')
// (18, 15, 'sp4_r_v_b_44')
// (18, 16, 'neigh_op_tnr_2')
// (18, 16, 'sp4_r_v_b_33')
// (18, 17, 'neigh_op_rgt_2')
// (18, 17, 'sp4_r_v_b_20')
// (18, 18, 'neigh_op_bnr_2')
// (18, 18, 'sp4_r_v_b_9')
// (19, 10, 'sp4_h_l_37')
// (19, 10, 'sp4_v_t_37')
// (19, 11, 'sp4_v_b_37')
// (19, 12, 'sp4_v_b_24')
// (19, 13, 'sp4_v_b_13')
// (19, 14, 'sp4_v_b_0')
// (19, 14, 'sp4_v_t_44')
// (19, 15, 'sp4_v_b_44')
// (19, 16, 'neigh_op_top_2')
// (19, 16, 'sp4_v_b_33')
// (19, 17, 'lutff_2/out')
// (19, 17, 'sp4_v_b_20')
// (19, 18, 'neigh_op_bot_2')
// (19, 18, 'sp4_v_b_9')
// (20, 16, 'neigh_op_tnl_2')
// (20, 17, 'neigh_op_lft_2')
// (20, 18, 'neigh_op_bnl_2')

reg n930 = 0;
// (15, 10, 'sp4_h_r_8')
// (16, 9, 'neigh_op_tnr_0')
// (16, 10, 'neigh_op_rgt_0')
// (16, 10, 'sp4_h_r_21')
// (16, 10, 'sp4_h_r_5')
// (16, 11, 'neigh_op_bnr_0')
// (16, 15, 'sp4_r_v_b_37')
// (16, 16, 'sp4_r_v_b_24')
// (16, 17, 'sp4_r_v_b_13')
// (16, 18, 'sp4_r_v_b_0')
// (16, 25, 'sp4_r_v_b_39')
// (16, 26, 'sp4_r_v_b_26')
// (16, 27, 'sp4_r_v_b_15')
// (16, 28, 'sp4_r_v_b_2')
// (17, 6, 'sp12_v_t_23')
// (17, 7, 'sp12_v_b_23')
// (17, 8, 'sp12_v_b_20')
// (17, 8, 'sp4_r_v_b_41')
// (17, 9, 'neigh_op_top_0')
// (17, 9, 'sp12_v_b_19')
// (17, 9, 'sp4_r_v_b_28')
// (17, 10, 'local_g0_0')
// (17, 10, 'lutff_0/in_0')
// (17, 10, 'lutff_0/out')
// (17, 10, 'sp12_v_b_16')
// (17, 10, 'sp4_h_r_16')
// (17, 10, 'sp4_h_r_32')
// (17, 10, 'sp4_r_v_b_17')
// (17, 11, 'local_g0_0')
// (17, 11, 'lutff_2/in_0')
// (17, 11, 'lutff_4/in_0')
// (17, 11, 'neigh_op_bot_0')
// (17, 11, 'sp12_v_b_15')
// (17, 11, 'sp4_r_v_b_4')
// (17, 12, 'sp12_v_b_12')
// (17, 12, 'sp4_r_v_b_41')
// (17, 12, 'sp4_r_v_b_42')
// (17, 13, 'local_g1_4')
// (17, 13, 'lutff_3/in_0')
// (17, 13, 'sp12_v_b_11')
// (17, 13, 'sp4_r_v_b_28')
// (17, 13, 'sp4_r_v_b_31')
// (17, 14, 'sp12_v_b_8')
// (17, 14, 'sp4_r_v_b_17')
// (17, 14, 'sp4_r_v_b_18')
// (17, 14, 'sp4_v_t_37')
// (17, 15, 'sp12_v_b_7')
// (17, 15, 'sp4_r_v_b_4')
// (17, 15, 'sp4_r_v_b_7')
// (17, 15, 'sp4_v_b_37')
// (17, 16, 'local_g2_5')
// (17, 16, 'lutff_5/in_0')
// (17, 16, 'sp12_v_b_4')
// (17, 16, 'sp4_r_v_b_37')
// (17, 16, 'sp4_v_b_24')
// (17, 17, 'local_g0_5')
// (17, 17, 'lutff_2/in_1')
// (17, 17, 'lutff_7/in_2')
// (17, 17, 'sp12_v_b_3')
// (17, 17, 'sp4_r_v_b_24')
// (17, 17, 'sp4_v_b_13')
// (17, 18, 'sp12_v_b_0')
// (17, 18, 'sp12_v_t_23')
// (17, 18, 'sp4_h_r_6')
// (17, 18, 'sp4_r_v_b_13')
// (17, 18, 'sp4_v_b_0')
// (17, 19, 'sp12_v_b_23')
// (17, 19, 'sp4_r_v_b_0')
// (17, 20, 'sp12_v_b_20')
// (17, 20, 'sp4_h_r_8')
// (17, 21, 'sp12_v_b_19')
// (17, 22, 'sp12_v_b_16')
// (17, 23, 'sp12_v_b_15')
// (17, 24, 'sp12_v_b_12')
// (17, 24, 'sp4_h_r_2')
// (17, 24, 'sp4_v_t_39')
// (17, 25, 'sp12_v_b_11')
// (17, 25, 'sp4_v_b_39')
// (17, 26, 'sp12_v_b_8')
// (17, 26, 'sp4_v_b_26')
// (17, 27, 'sp12_v_b_7')
// (17, 27, 'sp4_v_b_15')
// (17, 28, 'sp12_v_b_4')
// (17, 28, 'sp4_v_b_2')
// (17, 29, 'sp12_v_b_3')
// (17, 30, 'sp12_v_b_0')
// (18, 7, 'sp4_v_t_41')
// (18, 8, 'sp4_v_b_41')
// (18, 9, 'neigh_op_tnl_0')
// (18, 9, 'sp4_v_b_28')
// (18, 10, 'neigh_op_lft_0')
// (18, 10, 'sp4_h_r_29')
// (18, 10, 'sp4_h_r_45')
// (18, 10, 'sp4_v_b_17')
// (18, 11, 'neigh_op_bnl_0')
// (18, 11, 'sp4_r_v_b_39')
// (18, 11, 'sp4_v_b_4')
// (18, 11, 'sp4_v_t_41')
// (18, 11, 'sp4_v_t_42')
// (18, 12, 'sp4_r_v_b_26')
// (18, 12, 'sp4_v_b_41')
// (18, 12, 'sp4_v_b_42')
// (18, 13, 'local_g3_7')
// (18, 13, 'lutff_2/in_0')
// (18, 13, 'lutff_6/in_0')
// (18, 13, 'sp4_r_v_b_15')
// (18, 13, 'sp4_v_b_28')
// (18, 13, 'sp4_v_b_31')
// (18, 14, 'local_g0_1')
// (18, 14, 'local_g1_1')
// (18, 14, 'lutff_2/in_0')
// (18, 14, 'lutff_4/in_1')
// (18, 14, 'sp4_r_v_b_2')
// (18, 14, 'sp4_v_b_17')
// (18, 14, 'sp4_v_b_18')
// (18, 15, 'sp4_h_r_10')
// (18, 15, 'sp4_r_v_b_39')
// (18, 15, 'sp4_v_b_4')
// (18, 15, 'sp4_v_b_7')
// (18, 15, 'sp4_v_t_37')
// (18, 16, 'local_g3_5')
// (18, 16, 'lutff_0/in_2')
// (18, 16, 'sp4_r_v_b_26')
// (18, 16, 'sp4_v_b_37')
// (18, 17, 'local_g2_0')
// (18, 17, 'lutff_5/in_1')
// (18, 17, 'sp4_r_v_b_15')
// (18, 17, 'sp4_v_b_24')
// (18, 18, 'local_g0_3')
// (18, 18, 'lutff_6/in_1')
// (18, 18, 'sp4_h_r_19')
// (18, 18, 'sp4_r_v_b_2')
// (18, 18, 'sp4_v_b_13')
// (18, 19, 'sp4_h_r_6')
// (18, 19, 'sp4_v_b_0')
// (18, 20, 'local_g0_5')
// (18, 20, 'lutff_1/in_0')
// (18, 20, 'lutff_7/in_0')
// (18, 20, 'sp4_h_r_21')
// (18, 24, 'local_g0_7')
// (18, 24, 'local_g1_7')
// (18, 24, 'lutff_4/in_0')
// (18, 24, 'lutff_7/in_0')
// (18, 24, 'sp4_h_r_15')
// (19, 10, 'sp4_h_l_45')
// (19, 10, 'sp4_h_r_40')
// (19, 10, 'sp4_h_r_8')
// (19, 10, 'sp4_v_t_39')
// (19, 11, 'sp4_r_v_b_39')
// (19, 11, 'sp4_v_b_39')
// (19, 12, 'sp4_r_v_b_26')
// (19, 12, 'sp4_v_b_26')
// (19, 13, 'sp4_r_v_b_15')
// (19, 13, 'sp4_v_b_15')
// (19, 14, 'sp4_r_v_b_2')
// (19, 14, 'sp4_v_b_2')
// (19, 14, 'sp4_v_t_39')
// (19, 15, 'sp4_h_r_23')
// (19, 15, 'sp4_r_v_b_45')
// (19, 15, 'sp4_v_b_39')
// (19, 16, 'sp4_r_v_b_32')
// (19, 16, 'sp4_v_b_26')
// (19, 17, 'local_g0_7')
// (19, 17, 'local_g3_5')
// (19, 17, 'lutff_3/in_0')
// (19, 17, 'lutff_4/in_0')
// (19, 17, 'sp4_r_v_b_21')
// (19, 17, 'sp4_v_b_15')
// (19, 18, 'sp4_h_r_30')
// (19, 18, 'sp4_r_v_b_8')
// (19, 18, 'sp4_v_b_2')
// (19, 19, 'sp4_h_r_19')
// (19, 20, 'sp4_h_r_32')
// (19, 24, 'sp4_h_r_26')
// (20, 10, 'sp4_h_l_40')
// (20, 10, 'sp4_h_r_21')
// (20, 10, 'sp4_h_r_8')
// (20, 10, 'sp4_v_t_39')
// (20, 11, 'sp4_v_b_39')
// (20, 12, 'sp4_v_b_26')
// (20, 13, 'local_g0_7')
// (20, 13, 'lutff_2/in_1')
// (20, 13, 'lutff_4/in_1')
// (20, 13, 'sp4_v_b_15')
// (20, 14, 'local_g0_2')
// (20, 14, 'local_g1_2')
// (20, 14, 'lutff_3/in_0')
// (20, 14, 'lutff_6/in_0')
// (20, 14, 'sp4_h_r_2')
// (20, 14, 'sp4_v_b_2')
// (20, 14, 'sp4_v_t_45')
// (20, 15, 'sp4_h_r_34')
// (20, 15, 'sp4_v_b_45')
// (20, 16, 'sp4_v_b_32')
// (20, 17, 'sp4_v_b_21')
// (20, 18, 'sp4_h_r_43')
// (20, 18, 'sp4_v_b_8')
// (20, 19, 'sp4_h_r_30')
// (20, 20, 'sp4_h_r_45')
// (20, 21, 'sp4_r_v_b_39')
// (20, 22, 'sp4_r_v_b_26')
// (20, 23, 'sp4_r_v_b_15')
// (20, 24, 'sp4_h_r_39')
// (20, 24, 'sp4_r_v_b_2')
// (21, 10, 'sp4_h_r_21')
// (21, 10, 'sp4_h_r_32')
// (21, 14, 'sp4_h_r_15')
// (21, 15, 'local_g2_7')
// (21, 15, 'lutff_2/in_1')
// (21, 15, 'lutff_4/in_1')
// (21, 15, 'sp4_h_r_47')
// (21, 16, 'sp4_r_v_b_37')
// (21, 17, 'sp4_r_v_b_24')
// (21, 18, 'sp4_h_l_43')
// (21, 18, 'sp4_r_v_b_13')
// (21, 19, 'local_g1_0')
// (21, 19, 'local_g3_3')
// (21, 19, 'lutff_0/in_0')
// (21, 19, 'lutff_3/in_0')
// (21, 19, 'sp4_h_r_43')
// (21, 19, 'sp4_r_v_b_0')
// (21, 20, 'sp4_h_l_45')
// (21, 20, 'sp4_h_r_11')
// (21, 20, 'sp4_v_t_39')
// (21, 21, 'local_g2_7')
// (21, 21, 'lutff_1/in_0')
// (21, 21, 'lutff_7/in_0')
// (21, 21, 'sp4_v_b_39')
// (21, 22, 'sp4_v_b_26')
// (21, 23, 'sp4_v_b_15')
// (21, 24, 'sp4_h_l_39')
// (21, 24, 'sp4_v_b_2')
// (22, 10, 'sp4_h_r_32')
// (22, 10, 'sp4_h_r_45')
// (22, 11, 'sp4_r_v_b_36')
// (22, 12, 'sp4_r_v_b_25')
// (22, 13, 'sp4_r_v_b_12')
// (22, 14, 'sp4_h_r_26')
// (22, 14, 'sp4_r_v_b_1')
// (22, 15, 'sp4_h_l_47')
// (22, 15, 'sp4_r_v_b_36')
// (22, 15, 'sp4_r_v_b_41')
// (22, 15, 'sp4_v_t_37')
// (22, 16, 'sp4_r_v_b_25')
// (22, 16, 'sp4_r_v_b_28')
// (22, 16, 'sp4_v_b_37')
// (22, 17, 'local_g3_1')
// (22, 17, 'lutff_2/in_0')
// (22, 17, 'lutff_4/in_0')
// (22, 17, 'sp4_r_v_b_12')
// (22, 17, 'sp4_r_v_b_17')
// (22, 17, 'sp4_v_b_24')
// (22, 18, 'local_g1_1')
// (22, 18, 'local_g1_4')
// (22, 18, 'lutff_3/in_0')
// (22, 18, 'lutff_4/in_0')
// (22, 18, 'sp4_r_v_b_1')
// (22, 18, 'sp4_r_v_b_4')
// (22, 18, 'sp4_v_b_13')
// (22, 19, 'sp4_h_l_43')
// (22, 19, 'sp4_v_b_0')
// (22, 20, 'local_g0_6')
// (22, 20, 'lutff_3/in_1')
// (22, 20, 'sp4_h_r_22')
// (23, 10, 'sp4_h_l_45')
// (23, 10, 'sp4_h_r_45')
// (23, 10, 'sp4_v_t_36')
// (23, 11, 'sp4_v_b_36')
// (23, 12, 'sp4_v_b_25')
// (23, 13, 'sp4_v_b_12')
// (23, 14, 'sp4_h_r_39')
// (23, 14, 'sp4_v_b_1')
// (23, 14, 'sp4_v_t_36')
// (23, 14, 'sp4_v_t_41')
// (23, 15, 'sp4_v_b_36')
// (23, 15, 'sp4_v_b_41')
// (23, 16, 'sp4_v_b_25')
// (23, 16, 'sp4_v_b_28')
// (23, 17, 'sp4_v_b_12')
// (23, 17, 'sp4_v_b_17')
// (23, 18, 'sp4_v_b_1')
// (23, 18, 'sp4_v_b_4')
// (23, 20, 'sp4_h_r_35')
// (24, 10, 'sp4_h_l_45')
// (24, 14, 'sp4_h_l_39')
// (24, 20, 'sp4_h_r_46')
// (25, 20, 'sp4_h_l_46')

reg n931 = 0;
// (15, 11, 'local_g1_0')
// (15, 11, 'lutff_0/in_3')
// (15, 11, 'sp4_h_r_8')
// (16, 11, 'sp4_h_r_21')
// (17, 11, 'sp4_h_r_32')
// (18, 7, 'neigh_op_tnr_3')
// (18, 8, 'neigh_op_rgt_3')
// (18, 8, 'sp4_r_v_b_38')
// (18, 9, 'neigh_op_bnr_3')
// (18, 9, 'sp4_r_v_b_27')
// (18, 10, 'sp4_r_v_b_14')
// (18, 11, 'sp4_h_r_45')
// (18, 11, 'sp4_r_v_b_3')
// (19, 7, 'neigh_op_top_3')
// (19, 7, 'sp4_v_t_38')
// (19, 8, 'lutff_3/out')
// (19, 8, 'sp4_v_b_38')
// (19, 9, 'neigh_op_bot_3')
// (19, 9, 'sp4_v_b_27')
// (19, 10, 'sp4_v_b_14')
// (19, 11, 'sp4_h_l_45')
// (19, 11, 'sp4_v_b_3')
// (20, 7, 'neigh_op_tnl_3')
// (20, 8, 'neigh_op_lft_3')
// (20, 9, 'neigh_op_bnl_3')

wire n932;
// (15, 11, 'neigh_op_tnr_6')
// (15, 12, 'neigh_op_rgt_6')
// (15, 13, 'neigh_op_bnr_6')
// (16, 11, 'neigh_op_top_6')
// (16, 12, 'lutff_6/out')
// (16, 12, 'sp4_r_v_b_45')
// (16, 13, 'local_g1_6')
// (16, 13, 'lutff_0/in_1')
// (16, 13, 'lutff_5/in_2')
// (16, 13, 'neigh_op_bot_6')
// (16, 13, 'sp4_r_v_b_32')
// (16, 14, 'sp4_r_v_b_21')
// (16, 15, 'sp4_r_v_b_8')
// (17, 11, 'neigh_op_tnl_6')
// (17, 11, 'sp4_v_t_45')
// (17, 12, 'neigh_op_lft_6')
// (17, 12, 'sp4_v_b_45')
// (17, 13, 'neigh_op_bnl_6')
// (17, 13, 'sp4_v_b_32')
// (17, 14, 'sp4_v_b_21')
// (17, 15, 'sp4_h_r_8')
// (17, 15, 'sp4_v_b_8')
// (18, 15, 'sp4_h_r_21')
// (19, 15, 'sp4_h_r_32')
// (20, 15, 'local_g3_5')
// (20, 15, 'lutff_0/in_2')
// (20, 15, 'lutff_1/in_1')
// (20, 15, 'lutff_2/in_2')
// (20, 15, 'sp4_h_r_45')
// (21, 15, 'sp4_h_l_45')

wire n933;
// (15, 11, 'sp4_h_r_3')
// (16, 7, 'sp4_r_v_b_43')
// (16, 8, 'sp4_r_v_b_30')
// (16, 9, 'local_g3_3')
// (16, 9, 'lutff_global/cen')
// (16, 9, 'sp4_r_v_b_19')
// (16, 10, 'sp4_r_v_b_6')
// (16, 11, 'sp4_h_r_14')
// (17, 6, 'sp4_v_t_43')
// (17, 7, 'sp4_v_b_43')
// (17, 8, 'sp4_v_b_30')
// (17, 9, 'sp4_v_b_19')
// (17, 10, 'sp4_h_r_6')
// (17, 10, 'sp4_v_b_6')
// (17, 11, 'local_g3_3')
// (17, 11, 'lutff_global/cen')
// (17, 11, 'sp4_h_r_27')
// (18, 10, 'sp4_h_r_19')
// (18, 11, 'sp4_h_r_38')
// (18, 12, 'sp4_r_v_b_38')
// (18, 13, 'sp4_r_v_b_27')
// (18, 14, 'sp4_r_v_b_14')
// (18, 15, 'sp4_r_v_b_3')
// (19, 10, 'sp4_h_r_30')
// (19, 11, 'sp4_h_l_38')
// (19, 11, 'sp4_v_t_38')
// (19, 12, 'sp4_v_b_38')
// (19, 13, 'sp4_v_b_27')
// (19, 14, 'neigh_op_tnr_7')
// (19, 14, 'sp4_v_b_14')
// (19, 15, 'neigh_op_rgt_7')
// (19, 15, 'sp4_h_r_3')
// (19, 15, 'sp4_v_b_3')
// (19, 16, 'neigh_op_bnr_7')
// (20, 10, 'sp4_h_r_43')
// (20, 11, 'sp4_r_v_b_43')
// (20, 12, 'sp4_r_v_b_30')
// (20, 13, 'local_g3_3')
// (20, 13, 'lutff_global/cen')
// (20, 13, 'sp4_r_v_b_19')
// (20, 14, 'neigh_op_top_7')
// (20, 14, 'sp4_r_v_b_6')
// (20, 15, 'lutff_7/out')
// (20, 15, 'sp4_h_r_14')
// (20, 15, 'sp4_r_v_b_47')
// (20, 16, 'neigh_op_bot_7')
// (20, 16, 'sp4_r_v_b_34')
// (20, 17, 'sp4_r_v_b_23')
// (20, 18, 'sp4_r_v_b_10')
// (21, 10, 'sp4_h_l_43')
// (21, 10, 'sp4_v_t_43')
// (21, 11, 'sp4_v_b_43')
// (21, 12, 'sp4_v_b_30')
// (21, 13, 'sp4_v_b_19')
// (21, 14, 'neigh_op_tnl_7')
// (21, 14, 'sp4_v_b_6')
// (21, 14, 'sp4_v_t_47')
// (21, 15, 'local_g3_3')
// (21, 15, 'lutff_global/cen')
// (21, 15, 'neigh_op_lft_7')
// (21, 15, 'sp4_h_r_27')
// (21, 15, 'sp4_v_b_47')
// (21, 16, 'neigh_op_bnl_7')
// (21, 16, 'sp4_v_b_34')
// (21, 17, 'sp4_v_b_23')
// (21, 18, 'sp4_v_b_10')
// (22, 15, 'sp4_h_r_38')
// (23, 15, 'sp4_h_l_38')

wire n934;
// (15, 12, 'local_g3_4')
// (15, 12, 'lutff_1/in_0')
// (15, 12, 'sp4_r_v_b_44')
// (15, 13, 'sp4_r_v_b_33')
// (15, 14, 'sp4_r_v_b_20')
// (15, 15, 'sp4_r_v_b_9')
// (16, 11, 'sp4_v_t_44')
// (16, 12, 'sp4_v_b_44')
// (16, 13, 'sp4_v_b_33')
// (16, 14, 'sp4_v_b_20')
// (16, 15, 'sp4_h_r_9')
// (16, 15, 'sp4_v_b_9')
// (17, 15, 'sp4_h_r_20')
// (18, 15, 'sp4_h_r_33')
// (19, 15, 'sp4_h_r_44')
// (19, 16, 'sp4_r_v_b_44')
// (19, 17, 'neigh_op_tnr_2')
// (19, 17, 'sp4_r_v_b_33')
// (19, 18, 'neigh_op_rgt_2')
// (19, 18, 'sp4_r_v_b_20')
// (19, 19, 'neigh_op_bnr_2')
// (19, 19, 'sp4_r_v_b_9')
// (20, 15, 'sp4_h_l_44')
// (20, 15, 'sp4_v_t_44')
// (20, 16, 'sp4_v_b_44')
// (20, 17, 'neigh_op_top_2')
// (20, 17, 'sp4_v_b_33')
// (20, 18, 'lutff_2/out')
// (20, 18, 'sp4_v_b_20')
// (20, 19, 'neigh_op_bot_2')
// (20, 19, 'sp4_v_b_9')
// (21, 17, 'neigh_op_tnl_2')
// (21, 18, 'neigh_op_lft_2')
// (21, 19, 'neigh_op_bnl_2')

wire n935;
// (15, 12, 'neigh_op_tnr_2')
// (15, 13, 'neigh_op_rgt_2')
// (15, 13, 'sp4_r_v_b_36')
// (15, 14, 'local_g1_2')
// (15, 14, 'lutff_1/in_0')
// (15, 14, 'neigh_op_bnr_2')
// (15, 14, 'sp4_r_v_b_25')
// (15, 15, 'sp4_r_v_b_12')
// (15, 16, 'sp4_r_v_b_1')
// (16, 3, 'sp12_v_t_23')
// (16, 4, 'sp12_v_b_23')
// (16, 5, 'sp12_v_b_20')
// (16, 6, 'sp12_v_b_19')
// (16, 7, 'sp12_v_b_16')
// (16, 8, 'sp12_v_b_15')
// (16, 9, 'sp12_v_b_12')
// (16, 10, 'sp12_v_b_11')
// (16, 11, 'sp12_v_b_8')
// (16, 12, 'neigh_op_top_2')
// (16, 12, 'sp12_v_b_7')
// (16, 12, 'sp4_v_t_36')
// (16, 13, 'lutff_2/out')
// (16, 13, 'sp12_v_b_4')
// (16, 13, 'sp4_v_b_36')
// (16, 14, 'local_g3_1')
// (16, 14, 'lutff_0/in_2')
// (16, 14, 'lutff_1/in_1')
// (16, 14, 'neigh_op_bot_2')
// (16, 14, 'sp12_v_b_3')
// (16, 14, 'sp4_v_b_25')
// (16, 15, 'sp12_h_r_0')
// (16, 15, 'sp12_v_b_0')
// (16, 15, 'sp4_v_b_12')
// (16, 16, 'sp4_v_b_1')
// (17, 12, 'neigh_op_tnl_2')
// (17, 13, 'neigh_op_lft_2')
// (17, 14, 'neigh_op_bnl_2')
// (17, 15, 'sp12_h_r_3')
// (18, 15, 'local_g0_4')
// (18, 15, 'lutff_0/in_2')
// (18, 15, 'sp12_h_r_4')
// (19, 15, 'sp12_h_r_7')
// (20, 15, 'sp12_h_r_8')
// (21, 15, 'sp12_h_r_11')
// (22, 15, 'sp12_h_r_12')
// (23, 15, 'sp12_h_r_15')
// (24, 15, 'sp12_h_r_16')
// (25, 15, 'sp12_h_r_19')
// (26, 15, 'sp12_h_r_20')
// (27, 15, 'sp12_h_r_23')
// (28, 15, 'sp12_h_l_23')

wire n936;
// (15, 12, 'neigh_op_tnr_4')
// (15, 13, 'neigh_op_rgt_4')
// (15, 14, 'neigh_op_bnr_4')
// (16, 12, 'neigh_op_top_4')
// (16, 13, 'lutff_4/out')
// (16, 13, 'sp12_h_r_0')
// (16, 13, 'sp12_v_t_23')
// (16, 14, 'neigh_op_bot_4')
// (16, 14, 'sp12_v_b_23')
// (16, 15, 'sp12_v_b_20')
// (16, 16, 'sp12_v_b_19')
// (16, 17, 'sp12_v_b_16')
// (16, 18, 'sp12_v_b_15')
// (16, 19, 'sp12_v_b_12')
// (16, 20, 'local_g3_3')
// (16, 20, 'lutff_4/in_2')
// (16, 20, 'lutff_5/in_1')
// (16, 20, 'sp12_v_b_11')
// (16, 21, 'sp12_v_b_8')
// (16, 22, 'sp12_v_b_7')
// (16, 23, 'sp12_v_b_4')
// (16, 24, 'sp12_v_b_3')
// (16, 25, 'sp12_v_b_0')
// (17, 12, 'neigh_op_tnl_4')
// (17, 13, 'neigh_op_lft_4')
// (17, 13, 'sp12_h_r_3')
// (17, 14, 'neigh_op_bnl_4')
// (18, 13, 'sp12_h_r_4')
// (19, 13, 'sp12_h_r_7')
// (20, 13, 'sp12_h_r_8')
// (21, 13, 'sp12_h_r_11')
// (22, 13, 'sp12_h_r_12')
// (23, 13, 'sp12_h_r_15')
// (24, 13, 'sp12_h_r_16')
// (25, 13, 'sp12_h_r_19')
// (26, 13, 'sp12_h_r_20')
// (27, 13, 'sp12_h_r_23')
// (28, 13, 'sp12_h_l_23')

wire n937;
// (15, 12, 'neigh_op_tnr_6')
// (15, 13, 'local_g0_1')
// (15, 13, 'lutff_1/in_0')
// (15, 13, 'neigh_op_rgt_6')
// (15, 13, 'sp4_h_r_1')
// (15, 14, 'neigh_op_bnr_6')
// (16, 12, 'neigh_op_top_6')
// (16, 13, 'lutff_6/out')
// (16, 13, 'sp4_h_r_12')
// (16, 13, 'sp4_r_v_b_45')
// (16, 14, 'local_g1_6')
// (16, 14, 'lutff_4/in_1')
// (16, 14, 'neigh_op_bot_6')
// (16, 14, 'sp4_r_v_b_32')
// (16, 15, 'sp4_r_v_b_21')
// (16, 16, 'sp4_r_v_b_8')
// (16, 17, 'sp4_r_v_b_46')
// (16, 18, 'sp4_r_v_b_35')
// (16, 19, 'sp4_r_v_b_22')
// (16, 20, 'local_g2_3')
// (16, 20, 'lutff_2/in_3')
// (16, 20, 'lutff_3/in_0')
// (16, 20, 'sp4_r_v_b_11')
// (17, 12, 'neigh_op_tnl_6')
// (17, 12, 'sp4_v_t_45')
// (17, 13, 'neigh_op_lft_6')
// (17, 13, 'sp4_h_r_25')
// (17, 13, 'sp4_v_b_45')
// (17, 14, 'neigh_op_bnl_6')
// (17, 14, 'sp4_v_b_32')
// (17, 15, 'sp4_v_b_21')
// (17, 16, 'sp4_v_b_8')
// (17, 16, 'sp4_v_t_46')
// (17, 17, 'sp4_v_b_46')
// (17, 18, 'sp4_v_b_35')
// (17, 19, 'sp4_v_b_22')
// (17, 20, 'sp4_h_r_11')
// (17, 20, 'sp4_v_b_11')
// (18, 13, 'sp4_h_r_36')
// (18, 20, 'sp4_h_r_22')
// (19, 13, 'sp4_h_l_36')
// (19, 20, 'local_g3_3')
// (19, 20, 'lutff_7/in_3')
// (19, 20, 'sp4_h_r_35')
// (20, 20, 'sp4_h_r_46')
// (21, 20, 'sp4_h_l_46')

wire n938;
// (15, 12, 'neigh_op_tnr_7')
// (15, 12, 'sp4_r_v_b_43')
// (15, 13, 'neigh_op_rgt_7')
// (15, 13, 'sp4_r_v_b_30')
// (15, 14, 'neigh_op_bnr_7')
// (15, 14, 'sp4_r_v_b_19')
// (15, 15, 'sp4_r_v_b_6')
// (16, 8, 'sp12_v_t_22')
// (16, 9, 'sp12_v_b_22')
// (16, 10, 'sp12_v_b_21')
// (16, 11, 'local_g2_2')
// (16, 11, 'lutff_global/cen')
// (16, 11, 'sp12_v_b_18')
// (16, 11, 'sp4_h_r_11')
// (16, 11, 'sp4_v_t_43')
// (16, 12, 'neigh_op_top_7')
// (16, 12, 'sp12_v_b_17')
// (16, 12, 'sp4_v_b_43')
// (16, 13, 'lutff_7/out')
// (16, 13, 'sp12_v_b_14')
// (16, 13, 'sp4_v_b_30')
// (16, 14, 'neigh_op_bot_7')
// (16, 14, 'sp12_v_b_13')
// (16, 14, 'sp4_v_b_19')
// (16, 15, 'sp12_v_b_10')
// (16, 15, 'sp4_v_b_6')
// (16, 16, 'sp12_v_b_9')
// (16, 17, 'sp12_v_b_6')
// (16, 18, 'sp12_v_b_5')
// (16, 19, 'sp12_v_b_2')
// (16, 20, 'sp12_v_b_1')
// (17, 11, 'sp4_h_r_22')
// (17, 12, 'neigh_op_tnl_7')
// (17, 13, 'neigh_op_lft_7')
// (17, 14, 'neigh_op_bnl_7')
// (18, 11, 'sp4_h_r_35')
// (19, 11, 'sp4_h_r_46')
// (20, 11, 'sp4_h_l_46')
// (20, 11, 'sp4_h_r_7')
// (21, 11, 'sp4_h_r_18')
// (22, 11, 'sp4_h_r_31')
// (23, 11, 'local_g2_2')
// (23, 11, 'lutff_global/cen')
// (23, 11, 'sp4_h_r_42')
// (24, 11, 'sp4_h_l_42')

reg n939 = 0;
// (15, 12, 'sp4_h_r_2')
// (16, 12, 'sp4_h_r_15')
// (17, 12, 'local_g3_2')
// (17, 12, 'lutff_6/in_3')
// (17, 12, 'sp4_h_r_26')
// (18, 12, 'sp4_h_r_39')
// (19, 12, 'sp4_h_l_39')
// (19, 12, 'sp4_h_r_2')
// (20, 12, 'sp4_h_r_15')
// (21, 12, 'sp4_h_r_26')
// (22, 12, 'sp4_h_r_39')
// (22, 13, 'sp4_r_v_b_39')
// (22, 14, 'sp4_r_v_b_26')
// (22, 15, 'neigh_op_tnr_1')
// (22, 15, 'sp4_r_v_b_15')
// (22, 16, 'neigh_op_rgt_1')
// (22, 16, 'sp4_r_v_b_2')
// (22, 17, 'neigh_op_bnr_1')
// (23, 12, 'sp4_h_l_39')
// (23, 12, 'sp4_v_t_39')
// (23, 13, 'sp4_v_b_39')
// (23, 14, 'sp4_v_b_26')
// (23, 15, 'neigh_op_top_1')
// (23, 15, 'sp4_v_b_15')
// (23, 16, 'lutff_1/out')
// (23, 16, 'sp4_v_b_2')
// (23, 17, 'neigh_op_bot_1')
// (24, 15, 'neigh_op_tnl_1')
// (24, 16, 'neigh_op_lft_1')
// (24, 17, 'neigh_op_bnl_1')

reg n940 = 0;
// (15, 12, 'sp4_h_r_3')
// (16, 12, 'sp4_h_r_14')
// (17, 12, 'local_g2_3')
// (17, 12, 'lutff_4/in_3')
// (17, 12, 'sp4_h_r_27')
// (18, 9, 'sp4_r_v_b_38')
// (18, 10, 'neigh_op_tnr_7')
// (18, 10, 'sp4_r_v_b_27')
// (18, 11, 'neigh_op_rgt_7')
// (18, 11, 'sp4_r_v_b_14')
// (18, 12, 'neigh_op_bnr_7')
// (18, 12, 'sp4_h_r_38')
// (18, 12, 'sp4_r_v_b_3')
// (19, 8, 'sp4_v_t_38')
// (19, 9, 'sp4_v_b_38')
// (19, 10, 'neigh_op_top_7')
// (19, 10, 'sp4_v_b_27')
// (19, 11, 'lutff_7/out')
// (19, 11, 'sp4_v_b_14')
// (19, 12, 'neigh_op_bot_7')
// (19, 12, 'sp4_h_l_38')
// (19, 12, 'sp4_v_b_3')
// (20, 10, 'neigh_op_tnl_7')
// (20, 11, 'neigh_op_lft_7')
// (20, 12, 'neigh_op_bnl_7')

reg n941 = 0;
// (15, 12, 'sp4_h_r_4')
// (16, 12, 'sp4_h_r_17')
// (17, 12, 'local_g2_4')
// (17, 12, 'lutff_1/in_1')
// (17, 12, 'sp4_h_r_28')
// (18, 12, 'sp4_h_r_41')
// (19, 12, 'sp4_h_l_41')
// (19, 12, 'sp4_h_r_4')
// (20, 12, 'sp4_h_r_17')
// (21, 12, 'sp4_h_r_28')
// (22, 12, 'sp4_h_r_41')
// (22, 13, 'neigh_op_tnr_6')
// (22, 13, 'sp4_r_v_b_41')
// (22, 14, 'neigh_op_rgt_6')
// (22, 14, 'sp4_r_v_b_28')
// (22, 15, 'neigh_op_bnr_6')
// (22, 15, 'sp4_r_v_b_17')
// (22, 16, 'sp4_r_v_b_4')
// (23, 12, 'sp4_h_l_41')
// (23, 12, 'sp4_v_t_41')
// (23, 13, 'neigh_op_top_6')
// (23, 13, 'sp4_v_b_41')
// (23, 14, 'lutff_6/out')
// (23, 14, 'sp4_v_b_28')
// (23, 15, 'neigh_op_bot_6')
// (23, 15, 'sp4_v_b_17')
// (23, 16, 'sp4_v_b_4')
// (24, 13, 'neigh_op_tnl_6')
// (24, 14, 'neigh_op_lft_6')
// (24, 15, 'neigh_op_bnl_6')

reg n942 = 0;
// (15, 12, 'sp4_h_r_9')
// (16, 12, 'sp4_h_r_20')
// (17, 12, 'local_g3_1')
// (17, 12, 'lutff_1/in_3')
// (17, 12, 'sp4_h_r_33')
// (18, 12, 'sp4_h_r_44')
// (19, 12, 'sp4_h_l_44')
// (19, 12, 'sp4_h_r_1')
// (20, 12, 'sp4_h_r_12')
// (21, 12, 'sp4_h_r_25')
// (22, 12, 'sp4_h_r_36')
// (22, 13, 'sp4_r_v_b_36')
// (22, 14, 'neigh_op_tnr_6')
// (22, 14, 'sp4_r_v_b_25')
// (22, 15, 'neigh_op_rgt_6')
// (22, 15, 'sp4_r_v_b_12')
// (22, 16, 'neigh_op_bnr_6')
// (22, 16, 'sp4_r_v_b_1')
// (23, 12, 'sp4_h_l_36')
// (23, 12, 'sp4_v_t_36')
// (23, 13, 'sp4_v_b_36')
// (23, 14, 'neigh_op_top_6')
// (23, 14, 'sp4_v_b_25')
// (23, 15, 'lutff_6/out')
// (23, 15, 'sp4_v_b_12')
// (23, 16, 'neigh_op_bot_6')
// (23, 16, 'sp4_v_b_1')
// (24, 14, 'neigh_op_tnl_6')
// (24, 15, 'neigh_op_lft_6')
// (24, 16, 'neigh_op_bnl_6')

reg n943 = 0;
// (15, 12, 'sp4_r_v_b_46')
// (15, 13, 'local_g2_3')
// (15, 13, 'lutff_0/in_1')
// (15, 13, 'lutff_4/in_1')
// (15, 13, 'neigh_op_tnr_3')
// (15, 13, 'sp4_r_v_b_35')
// (15, 14, 'neigh_op_rgt_3')
// (15, 14, 'sp4_r_v_b_22')
// (15, 15, 'neigh_op_bnr_3')
// (15, 15, 'sp4_r_v_b_11')
// (16, 11, 'sp4_r_v_b_42')
// (16, 11, 'sp4_v_t_46')
// (16, 12, 'local_g0_7')
// (16, 12, 'lutff_2/in_1')
// (16, 12, 'sp4_r_v_b_31')
// (16, 12, 'sp4_v_b_46')
// (16, 13, 'neigh_op_top_3')
// (16, 13, 'sp4_r_v_b_18')
// (16, 13, 'sp4_v_b_35')
// (16, 14, 'local_g0_3')
// (16, 14, 'lutff_0/in_1')
// (16, 14, 'lutff_1/in_0')
// (16, 14, 'lutff_3/out')
// (16, 14, 'lutff_5/in_0')
// (16, 14, 'sp4_r_v_b_7')
// (16, 14, 'sp4_v_b_22')
// (16, 15, 'local_g1_3')
// (16, 15, 'lutff_0/in_2')
// (16, 15, 'lutff_3/in_1')
// (16, 15, 'neigh_op_bot_3')
// (16, 15, 'sp4_h_r_5')
// (16, 15, 'sp4_v_b_11')
// (17, 10, 'sp4_v_t_42')
// (17, 11, 'sp4_v_b_42')
// (17, 12, 'sp4_v_b_31')
// (17, 13, 'neigh_op_tnl_3')
// (17, 13, 'sp4_v_b_18')
// (17, 14, 'neigh_op_lft_3')
// (17, 14, 'sp4_v_b_7')
// (17, 15, 'neigh_op_bnl_3')
// (17, 15, 'sp4_h_r_16')
// (18, 15, 'local_g3_5')
// (18, 15, 'lutff_0/in_0')
// (18, 15, 'sp4_h_r_29')
// (19, 15, 'sp4_h_r_40')
// (20, 15, 'sp4_h_l_40')

wire n944;
// (15, 12, 'sp4_r_v_b_47')
// (15, 13, 'sp4_r_v_b_34')
// (15, 14, 'neigh_op_tnr_5')
// (15, 14, 'sp4_r_v_b_23')
// (15, 15, 'local_g2_2')
// (15, 15, 'lutff_global/cen')
// (15, 15, 'neigh_op_rgt_5')
// (15, 15, 'sp4_r_v_b_10')
// (15, 16, 'neigh_op_bnr_5')
// (16, 11, 'sp4_v_t_47')
// (16, 12, 'sp4_v_b_47')
// (16, 13, 'sp4_v_b_34')
// (16, 14, 'neigh_op_top_5')
// (16, 14, 'sp4_v_b_23')
// (16, 15, 'lutff_5/out')
// (16, 15, 'sp4_v_b_10')
// (16, 16, 'neigh_op_bot_5')
// (17, 14, 'neigh_op_tnl_5')
// (17, 15, 'neigh_op_lft_5')
// (17, 16, 'neigh_op_bnl_5')

wire n945;
// (15, 13, 'lutff_0/lout')
// (15, 13, 'lutff_1/in_2')

wire n946;
// (15, 13, 'lutff_1/lout')
// (15, 13, 'lutff_2/in_2')

wire n947;
// (15, 13, 'lutff_4/lout')
// (15, 13, 'lutff_5/in_2')

wire n948;
// (15, 13, 'neigh_op_tnr_5')
// (15, 13, 'sp4_r_v_b_39')
// (15, 14, 'neigh_op_rgt_5')
// (15, 14, 'sp4_r_v_b_26')
// (15, 15, 'neigh_op_bnr_5')
// (15, 15, 'sp4_r_v_b_15')
// (15, 16, 'sp4_r_v_b_2')
// (16, 12, 'sp4_h_r_2')
// (16, 12, 'sp4_v_t_39')
// (16, 13, 'neigh_op_top_5')
// (16, 13, 'sp4_v_b_39')
// (16, 14, 'local_g2_5')
// (16, 14, 'lutff_2/in_3')
// (16, 14, 'lutff_4/in_3')
// (16, 14, 'lutff_5/out')
// (16, 14, 'lutff_7/in_0')
// (16, 14, 'sp4_v_b_26')
// (16, 15, 'local_g1_5')
// (16, 15, 'lutff_2/in_0')
// (16, 15, 'lutff_5/in_3')
// (16, 15, 'neigh_op_bot_5')
// (16, 15, 'sp4_v_b_15')
// (16, 16, 'sp4_v_b_2')
// (17, 12, 'sp4_h_r_15')
// (17, 13, 'neigh_op_tnl_5')
// (17, 14, 'neigh_op_lft_5')
// (17, 15, 'neigh_op_bnl_5')
// (18, 12, 'sp4_h_r_26')
// (19, 12, 'local_g2_7')
// (19, 12, 'lutff_0/in_3')
// (19, 12, 'lutff_5/in_0')
// (19, 12, 'sp4_h_r_39')
// (19, 13, 'sp4_r_v_b_42')
// (19, 14, 'sp4_r_v_b_31')
// (19, 15, 'sp4_r_v_b_18')
// (19, 16, 'sp4_r_v_b_7')
// (20, 12, 'sp4_h_l_39')
// (20, 12, 'sp4_v_t_42')
// (20, 13, 'sp4_v_b_42')
// (20, 14, 'sp4_v_b_31')
// (20, 15, 'local_g1_2')
// (20, 15, 'lutff_2/in_3')
// (20, 15, 'sp4_v_b_18')
// (20, 16, 'sp4_v_b_7')

wire n949;
// (15, 13, 'neigh_op_tnr_7')
// (15, 13, 'sp4_r_v_b_43')
// (15, 14, 'neigh_op_rgt_7')
// (15, 14, 'sp4_r_v_b_30')
// (15, 15, 'neigh_op_bnr_7')
// (15, 15, 'sp4_r_v_b_19')
// (15, 16, 'sp4_r_v_b_6')
// (16, 12, 'sp4_v_t_43')
// (16, 13, 'neigh_op_top_7')
// (16, 13, 'sp4_v_b_43')
// (16, 14, 'lutff_7/out')
// (16, 14, 'sp4_v_b_30')
// (16, 15, 'neigh_op_bot_7')
// (16, 15, 'sp4_v_b_19')
// (16, 16, 'sp4_h_r_6')
// (16, 16, 'sp4_v_b_6')
// (17, 13, 'neigh_op_tnl_7')
// (17, 14, 'neigh_op_lft_7')
// (17, 15, 'neigh_op_bnl_7')
// (17, 16, 'sp4_h_r_19')
// (18, 16, 'sp4_h_r_30')
// (19, 16, 'local_g3_3')
// (19, 16, 'lutff_global/cen')
// (19, 16, 'sp4_h_r_43')
// (20, 16, 'sp4_h_l_43')

wire n950;
// (15, 13, 'sp12_h_r_0')
// (16, 13, 'sp12_h_r_3')
// (17, 13, 'sp12_h_r_4')
// (18, 13, 'local_g0_7')
// (18, 13, 'lutff_2/in_1')
// (18, 13, 'sp12_h_r_7')
// (19, 13, 'sp12_h_r_8')
// (20, 13, 'sp12_h_r_11')
// (21, 13, 'sp12_h_r_12')
// (22, 12, 'neigh_op_tnr_4')
// (22, 13, 'neigh_op_rgt_4')
// (22, 13, 'sp12_h_r_15')
// (22, 14, 'neigh_op_bnr_4')
// (23, 12, 'neigh_op_top_4')
// (23, 13, 'lutff_4/out')
// (23, 13, 'sp12_h_r_16')
// (23, 14, 'neigh_op_bot_4')
// (24, 12, 'neigh_op_tnl_4')
// (24, 13, 'neigh_op_lft_4')
// (24, 13, 'sp12_h_r_19')
// (24, 14, 'neigh_op_bnl_4')
// (25, 13, 'sp12_h_r_20')
// (26, 13, 'sp12_h_r_23')
// (27, 13, 'sp12_h_l_23')

reg n951 = 0;
// (15, 13, 'sp4_h_r_11')
// (16, 13, 'sp4_h_r_22')
// (17, 13, 'local_g3_3')
// (17, 13, 'lutff_5/in_1')
// (17, 13, 'sp4_h_r_35')
// (18, 9, 'neigh_op_tnr_7')
// (18, 10, 'neigh_op_rgt_7')
// (18, 10, 'sp4_r_v_b_46')
// (18, 11, 'neigh_op_bnr_7')
// (18, 11, 'sp4_r_v_b_35')
// (18, 12, 'sp4_r_v_b_22')
// (18, 13, 'sp4_h_r_46')
// (18, 13, 'sp4_r_v_b_11')
// (19, 9, 'neigh_op_top_7')
// (19, 9, 'sp4_v_t_46')
// (19, 10, 'lutff_7/out')
// (19, 10, 'sp4_v_b_46')
// (19, 11, 'neigh_op_bot_7')
// (19, 11, 'sp4_v_b_35')
// (19, 12, 'sp4_v_b_22')
// (19, 13, 'sp4_h_l_46')
// (19, 13, 'sp4_v_b_11')
// (20, 9, 'neigh_op_tnl_7')
// (20, 10, 'neigh_op_lft_7')
// (20, 11, 'neigh_op_bnl_7')

reg n952 = 0;
// (15, 13, 'sp4_h_r_3')
// (16, 13, 'sp4_h_r_14')
// (17, 13, 'local_g2_3')
// (17, 13, 'lutff_6/in_3')
// (17, 13, 'sp4_h_r_27')
// (18, 13, 'sp4_h_r_38')
// (18, 14, 'sp4_r_v_b_38')
// (18, 15, 'neigh_op_tnr_7')
// (18, 15, 'sp4_r_v_b_27')
// (18, 16, 'neigh_op_rgt_7')
// (18, 16, 'sp4_r_v_b_14')
// (18, 17, 'neigh_op_bnr_7')
// (18, 17, 'sp4_r_v_b_3')
// (19, 13, 'sp4_h_l_38')
// (19, 13, 'sp4_v_t_38')
// (19, 14, 'sp4_v_b_38')
// (19, 15, 'neigh_op_top_7')
// (19, 15, 'sp4_v_b_27')
// (19, 16, 'lutff_7/out')
// (19, 16, 'sp4_v_b_14')
// (19, 17, 'neigh_op_bot_7')
// (19, 17, 'sp4_v_b_3')
// (20, 15, 'neigh_op_tnl_7')
// (20, 16, 'neigh_op_lft_7')
// (20, 17, 'neigh_op_bnl_7')

reg n953 = 0;
// (15, 13, 'sp4_h_r_4')
// (16, 13, 'sp4_h_r_17')
// (17, 13, 'sp4_h_r_28')
// (18, 13, 'local_g3_1')
// (18, 13, 'lutff_1/in_1')
// (18, 13, 'sp4_h_r_41')
// (19, 13, 'sp4_h_l_41')
// (19, 13, 'sp4_h_r_1')
// (20, 13, 'sp4_h_r_12')
// (21, 13, 'sp4_h_r_25')
// (22, 10, 'sp4_r_v_b_36')
// (22, 11, 'neigh_op_tnr_6')
// (22, 11, 'sp4_r_v_b_25')
// (22, 12, 'neigh_op_rgt_6')
// (22, 12, 'sp4_r_v_b_12')
// (22, 13, 'neigh_op_bnr_6')
// (22, 13, 'sp4_h_r_36')
// (22, 13, 'sp4_r_v_b_1')
// (23, 9, 'sp4_v_t_36')
// (23, 10, 'sp4_v_b_36')
// (23, 11, 'neigh_op_top_6')
// (23, 11, 'sp4_v_b_25')
// (23, 12, 'lutff_6/out')
// (23, 12, 'sp4_v_b_12')
// (23, 13, 'neigh_op_bot_6')
// (23, 13, 'sp4_h_l_36')
// (23, 13, 'sp4_v_b_1')
// (24, 11, 'neigh_op_tnl_6')
// (24, 12, 'neigh_op_lft_6')
// (24, 13, 'neigh_op_bnl_6')

reg n954 = 0;
// (15, 13, 'sp4_h_r_9')
// (16, 13, 'sp4_h_r_20')
// (17, 13, 'local_g3_1')
// (17, 13, 'lutff_1/in_1')
// (17, 13, 'sp4_h_r_33')
// (18, 9, 'neigh_op_tnr_6')
// (18, 10, 'neigh_op_rgt_6')
// (18, 10, 'sp4_r_v_b_44')
// (18, 11, 'neigh_op_bnr_6')
// (18, 11, 'sp4_r_v_b_33')
// (18, 12, 'sp4_r_v_b_20')
// (18, 13, 'sp4_h_r_44')
// (18, 13, 'sp4_r_v_b_9')
// (19, 9, 'neigh_op_top_6')
// (19, 9, 'sp4_v_t_44')
// (19, 10, 'lutff_6/out')
// (19, 10, 'sp4_v_b_44')
// (19, 11, 'neigh_op_bot_6')
// (19, 11, 'sp4_v_b_33')
// (19, 12, 'sp4_v_b_20')
// (19, 13, 'sp4_h_l_44')
// (19, 13, 'sp4_v_b_9')
// (20, 9, 'neigh_op_tnl_6')
// (20, 10, 'neigh_op_lft_6')
// (20, 11, 'neigh_op_bnl_6')

wire n955;
// (15, 14, 'lutff_0/lout')
// (15, 14, 'lutff_1/in_2')

wire n956;
// (15, 14, 'lutff_1/lout')
// (15, 14, 'lutff_2/in_2')

wire n957;
// (15, 14, 'lutff_6/lout')
// (15, 14, 'lutff_7/in_2')

wire n958;
// (15, 14, 'neigh_op_tnr_1')
// (15, 15, 'neigh_op_rgt_1')
// (15, 16, 'neigh_op_bnr_1')
// (16, 12, 'sp4_r_v_b_38')
// (16, 12, 'sp4_r_v_b_42')
// (16, 13, 'sp4_r_v_b_27')
// (16, 13, 'sp4_r_v_b_31')
// (16, 14, 'neigh_op_top_1')
// (16, 14, 'sp4_r_v_b_14')
// (16, 14, 'sp4_r_v_b_18')
// (16, 15, 'lutff_1/out')
// (16, 15, 'sp4_r_v_b_3')
// (16, 15, 'sp4_r_v_b_7')
// (16, 16, 'neigh_op_bot_1')
// (16, 16, 'sp4_r_v_b_46')
// (16, 17, 'sp4_r_v_b_35')
// (16, 18, 'sp4_r_v_b_22')
// (16, 19, 'sp4_r_v_b_11')
// (17, 11, 'sp4_v_t_38')
// (17, 11, 'sp4_v_t_42')
// (17, 12, 'sp4_v_b_38')
// (17, 12, 'sp4_v_b_42')
// (17, 13, 'sp4_v_b_27')
// (17, 13, 'sp4_v_b_31')
// (17, 14, 'local_g0_2')
// (17, 14, 'lutff_global/cen')
// (17, 14, 'neigh_op_tnl_1')
// (17, 14, 'sp4_v_b_14')
// (17, 14, 'sp4_v_b_18')
// (17, 15, 'neigh_op_lft_1')
// (17, 15, 'sp4_h_r_11')
// (17, 15, 'sp4_v_b_3')
// (17, 15, 'sp4_v_b_7')
// (17, 15, 'sp4_v_t_46')
// (17, 16, 'neigh_op_bnl_1')
// (17, 16, 'sp4_v_b_46')
// (17, 17, 'sp4_v_b_35')
// (17, 18, 'sp4_v_b_22')
// (17, 19, 'sp4_v_b_11')
// (18, 15, 'sp4_h_r_22')
// (19, 15, 'sp4_h_r_35')
// (20, 15, 'sp4_h_r_46')
// (20, 16, 'sp4_r_v_b_42')
// (20, 17, 'sp4_r_v_b_31')
// (20, 18, 'sp4_r_v_b_18')
// (20, 19, 'sp4_r_v_b_7')
// (21, 15, 'sp4_h_l_46')
// (21, 15, 'sp4_h_r_7')
// (21, 15, 'sp4_v_t_42')
// (21, 16, 'sp4_v_b_42')
// (21, 17, 'sp4_v_b_31')
// (21, 18, 'local_g0_2')
// (21, 18, 'lutff_global/cen')
// (21, 18, 'sp4_v_b_18')
// (21, 19, 'sp4_v_b_7')
// (22, 15, 'sp4_h_r_18')
// (23, 15, 'sp4_h_r_31')
// (24, 15, 'local_g2_2')
// (24, 15, 'lutff_global/cen')
// (24, 15, 'sp4_h_r_42')
// (25, 15, 'sp4_h_l_42')

wire n959;
// (15, 14, 'sp4_h_r_10')
// (16, 13, 'neigh_op_tnr_1')
// (16, 14, 'neigh_op_rgt_1')
// (16, 14, 'sp4_h_r_23')
// (16, 15, 'neigh_op_bnr_1')
// (17, 13, 'neigh_op_top_1')
// (17, 14, 'lutff_1/out')
// (17, 14, 'sp4_h_r_34')
// (17, 15, 'neigh_op_bot_1')
// (18, 13, 'neigh_op_tnl_1')
// (18, 14, 'neigh_op_lft_1')
// (18, 14, 'sp4_h_r_47')
// (18, 15, 'neigh_op_bnl_1')
// (18, 15, 'sp4_r_v_b_47')
// (18, 16, 'sp4_r_v_b_34')
// (18, 17, 'sp4_r_v_b_23')
// (18, 18, 'sp4_r_v_b_10')
// (19, 14, 'sp4_h_l_47')
// (19, 14, 'sp4_v_t_47')
// (19, 15, 'sp4_v_b_47')
// (19, 16, 'sp4_v_b_34')
// (19, 17, 'local_g1_7')
// (19, 17, 'lutff_0/in_0')
// (19, 17, 'sp4_v_b_23')
// (19, 18, 'sp4_v_b_10')

reg n960 = 0;
// (15, 14, 'sp4_h_r_4')
// (16, 14, 'sp4_h_r_17')
// (17, 14, 'sp4_h_r_28')
// (18, 14, 'local_g3_1')
// (18, 14, 'lutff_6/in_0')
// (18, 14, 'sp4_h_r_41')
// (19, 14, 'sp4_h_l_41')
// (19, 14, 'sp4_h_r_8')
// (20, 14, 'sp4_h_r_21')
// (21, 14, 'sp4_h_r_32')
// (22, 11, 'neigh_op_tnr_0')
// (22, 11, 'sp4_r_v_b_45')
// (22, 12, 'neigh_op_rgt_0')
// (22, 12, 'sp4_r_v_b_32')
// (22, 13, 'neigh_op_bnr_0')
// (22, 13, 'sp4_r_v_b_21')
// (22, 14, 'sp4_h_r_45')
// (22, 14, 'sp4_r_v_b_8')
// (23, 10, 'sp4_v_t_45')
// (23, 11, 'neigh_op_top_0')
// (23, 11, 'sp4_v_b_45')
// (23, 12, 'lutff_0/out')
// (23, 12, 'sp4_v_b_32')
// (23, 13, 'neigh_op_bot_0')
// (23, 13, 'sp4_v_b_21')
// (23, 14, 'sp4_h_l_45')
// (23, 14, 'sp4_v_b_8')
// (24, 11, 'neigh_op_tnl_0')
// (24, 12, 'neigh_op_lft_0')
// (24, 13, 'neigh_op_bnl_0')

reg n961 = 0;
// (15, 14, 'sp4_h_r_5')
// (16, 14, 'sp4_h_r_16')
// (17, 14, 'local_g3_5')
// (17, 14, 'lutff_1/in_3')
// (17, 14, 'sp4_h_r_29')
// (18, 14, 'sp4_h_r_40')
// (18, 15, 'sp4_r_v_b_40')
// (18, 16, 'sp4_r_v_b_29')
// (18, 17, 'sp4_r_v_b_16')
// (18, 18, 'neigh_op_tnr_4')
// (18, 18, 'sp4_r_v_b_5')
// (18, 19, 'neigh_op_rgt_4')
// (18, 19, 'sp4_r_v_b_40')
// (18, 20, 'neigh_op_bnr_4')
// (18, 20, 'sp4_r_v_b_29')
// (18, 21, 'sp4_r_v_b_16')
// (18, 22, 'sp4_r_v_b_5')
// (19, 14, 'sp4_h_l_40')
// (19, 14, 'sp4_v_t_40')
// (19, 15, 'sp4_v_b_40')
// (19, 16, 'sp4_v_b_29')
// (19, 17, 'sp4_v_b_16')
// (19, 18, 'neigh_op_top_4')
// (19, 18, 'sp4_v_b_5')
// (19, 18, 'sp4_v_t_40')
// (19, 19, 'lutff_4/out')
// (19, 19, 'sp4_v_b_40')
// (19, 20, 'neigh_op_bot_4')
// (19, 20, 'sp4_v_b_29')
// (19, 21, 'sp4_v_b_16')
// (19, 22, 'sp4_v_b_5')
// (20, 18, 'neigh_op_tnl_4')
// (20, 19, 'neigh_op_lft_4')
// (20, 20, 'neigh_op_bnl_4')

reg n962 = 0;
// (15, 14, 'sp4_r_v_b_44')
// (15, 15, 'neigh_op_tnr_2')
// (15, 15, 'sp4_r_v_b_33')
// (15, 16, 'neigh_op_rgt_2')
// (15, 16, 'sp4_r_v_b_20')
// (15, 17, 'neigh_op_bnr_2')
// (15, 17, 'sp4_r_v_b_9')
// (16, 13, 'sp4_h_r_2')
// (16, 13, 'sp4_v_t_44')
// (16, 14, 'sp4_v_b_44')
// (16, 15, 'neigh_op_top_2')
// (16, 15, 'sp4_v_b_33')
// (16, 16, 'lutff_2/out')
// (16, 16, 'sp4_v_b_20')
// (16, 17, 'neigh_op_bot_2')
// (16, 17, 'sp4_v_b_9')
// (17, 13, 'sp4_h_r_15')
// (17, 15, 'neigh_op_tnl_2')
// (17, 16, 'neigh_op_lft_2')
// (17, 17, 'neigh_op_bnl_2')
// (18, 13, 'sp4_h_r_26')
// (19, 13, 'sp4_h_r_39')
// (20, 13, 'sp4_h_l_39')
// (20, 13, 'sp4_h_r_2')
// (21, 13, 'local_g0_7')
// (21, 13, 'lutff_6/in_3')
// (21, 13, 'sp4_h_r_15')
// (22, 13, 'sp4_h_r_26')
// (23, 13, 'sp4_h_r_39')
// (24, 13, 'sp4_h_l_39')

reg n963 = 0;
// (15, 15, 'neigh_op_tnr_1')
// (15, 16, 'neigh_op_rgt_1')
// (15, 17, 'neigh_op_bnr_1')
// (16, 14, 'sp4_r_v_b_43')
// (16, 15, 'neigh_op_top_1')
// (16, 15, 'sp4_r_v_b_30')
// (16, 16, 'lutff_1/out')
// (16, 16, 'sp4_r_v_b_19')
// (16, 17, 'neigh_op_bot_1')
// (16, 17, 'sp4_r_v_b_6')
// (17, 13, 'sp4_h_r_6')
// (17, 13, 'sp4_v_t_43')
// (17, 14, 'sp4_v_b_43')
// (17, 15, 'neigh_op_tnl_1')
// (17, 15, 'sp4_v_b_30')
// (17, 16, 'neigh_op_lft_1')
// (17, 16, 'sp4_v_b_19')
// (17, 17, 'neigh_op_bnl_1')
// (17, 17, 'sp4_v_b_6')
// (18, 13, 'sp4_h_r_19')
// (19, 13, 'local_g3_6')
// (19, 13, 'lutff_2/in_3')
// (19, 13, 'sp4_h_r_30')
// (20, 13, 'sp4_h_r_43')
// (21, 13, 'sp4_h_l_43')

reg n964 = 0;
// (15, 15, 'neigh_op_tnr_3')
// (15, 16, 'neigh_op_rgt_3')
// (15, 16, 'sp4_h_r_11')
// (15, 17, 'neigh_op_bnr_3')
// (16, 15, 'neigh_op_top_3')
// (16, 16, 'lutff_3/out')
// (16, 16, 'sp4_h_r_22')
// (16, 17, 'neigh_op_bot_3')
// (17, 15, 'neigh_op_tnl_3')
// (17, 16, 'neigh_op_lft_3')
// (17, 16, 'sp4_h_r_35')
// (17, 17, 'neigh_op_bnl_3')
// (18, 16, 'sp4_h_r_46')
// (19, 16, 'sp4_h_l_46')
// (19, 16, 'sp4_h_r_7')
// (20, 16, 'sp4_h_r_18')
// (21, 16, 'local_g2_7')
// (21, 16, 'lutff_4/in_3')
// (21, 16, 'sp4_h_r_31')
// (22, 16, 'sp4_h_r_42')
// (23, 16, 'sp4_h_l_42')

reg n965 = 0;
// (15, 15, 'neigh_op_tnr_4')
// (15, 16, 'neigh_op_rgt_4')
// (15, 17, 'neigh_op_bnr_4')
// (16, 15, 'neigh_op_top_4')
// (16, 16, 'lutff_4/out')
// (16, 16, 'sp12_h_r_0')
// (16, 17, 'neigh_op_bot_4')
// (17, 15, 'neigh_op_tnl_4')
// (17, 16, 'neigh_op_lft_4')
// (17, 16, 'sp12_h_r_3')
// (17, 17, 'neigh_op_bnl_4')
// (18, 16, 'sp12_h_r_4')
// (19, 16, 'sp12_h_r_7')
// (20, 16, 'sp12_h_r_8')
// (21, 16, 'sp12_h_r_11')
// (22, 16, 'local_g1_4')
// (22, 16, 'lutff_6/in_3')
// (22, 16, 'sp12_h_r_12')
// (23, 16, 'sp12_h_r_15')
// (24, 16, 'sp12_h_r_16')
// (25, 16, 'sp12_h_r_19')
// (26, 16, 'sp12_h_r_20')
// (27, 16, 'sp12_h_r_23')
// (28, 16, 'sp12_h_l_23')

reg n966 = 0;
// (15, 15, 'neigh_op_tnr_5')
// (15, 16, 'neigh_op_rgt_5')
// (15, 17, 'neigh_op_bnr_5')
// (16, 15, 'neigh_op_top_5')
// (16, 15, 'sp4_r_v_b_38')
// (16, 16, 'lutff_5/out')
// (16, 16, 'sp4_r_v_b_27')
// (16, 17, 'neigh_op_bot_5')
// (16, 17, 'sp4_r_v_b_14')
// (16, 18, 'sp4_r_v_b_3')
// (17, 14, 'sp4_v_t_38')
// (17, 15, 'neigh_op_tnl_5')
// (17, 15, 'sp4_v_b_38')
// (17, 16, 'neigh_op_lft_5')
// (17, 16, 'sp4_v_b_27')
// (17, 17, 'neigh_op_bnl_5')
// (17, 17, 'sp4_v_b_14')
// (17, 18, 'sp4_h_r_9')
// (17, 18, 'sp4_v_b_3')
// (18, 18, 'sp4_h_r_20')
// (19, 18, 'local_g2_1')
// (19, 18, 'lutff_4/in_3')
// (19, 18, 'sp4_h_r_33')
// (20, 18, 'sp4_h_r_44')
// (21, 18, 'sp4_h_l_44')

reg n967 = 0;
// (15, 15, 'neigh_op_tnr_6')
// (15, 16, 'neigh_op_rgt_6')
// (15, 16, 'sp4_h_r_1')
// (15, 17, 'neigh_op_bnr_6')
// (16, 15, 'neigh_op_top_6')
// (16, 16, 'lutff_6/out')
// (16, 16, 'sp4_h_r_12')
// (16, 17, 'neigh_op_bot_6')
// (17, 15, 'neigh_op_tnl_6')
// (17, 16, 'neigh_op_lft_6')
// (17, 16, 'sp4_h_r_25')
// (17, 17, 'neigh_op_bnl_6')
// (18, 13, 'sp4_r_v_b_36')
// (18, 14, 'sp4_r_v_b_25')
// (18, 15, 'sp4_r_v_b_12')
// (18, 16, 'sp4_h_r_36')
// (18, 16, 'sp4_r_v_b_1')
// (19, 12, 'sp4_v_t_36')
// (19, 13, 'sp4_v_b_36')
// (19, 14, 'local_g2_1')
// (19, 14, 'lutff_4/in_3')
// (19, 14, 'sp4_v_b_25')
// (19, 15, 'sp4_v_b_12')
// (19, 16, 'sp4_h_l_36')
// (19, 16, 'sp4_v_b_1')

reg n968 = 0;
// (15, 15, 'neigh_op_tnr_7')
// (15, 16, 'neigh_op_rgt_7')
// (15, 17, 'neigh_op_bnr_7')
// (16, 14, 'sp4_r_v_b_39')
// (16, 15, 'neigh_op_top_7')
// (16, 15, 'sp4_r_v_b_26')
// (16, 16, 'lutff_7/out')
// (16, 16, 'sp4_r_v_b_15')
// (16, 17, 'neigh_op_bot_7')
// (16, 17, 'sp4_r_v_b_2')
// (17, 13, 'sp4_v_t_39')
// (17, 14, 'local_g3_7')
// (17, 14, 'lutff_7/in_3')
// (17, 14, 'sp4_v_b_39')
// (17, 15, 'neigh_op_tnl_7')
// (17, 15, 'sp4_v_b_26')
// (17, 16, 'neigh_op_lft_7')
// (17, 16, 'sp4_v_b_15')
// (17, 17, 'neigh_op_bnl_7')
// (17, 17, 'sp4_v_b_2')

reg n969 = 0;
// (15, 15, 'sp4_h_r_6')
// (16, 15, 'sp4_h_r_19')
// (17, 15, 'local_g3_6')
// (17, 15, 'lutff_6/in_3')
// (17, 15, 'sp4_h_r_30')
// (18, 15, 'sp4_h_r_43')
// (18, 16, 'sp4_r_v_b_37')
// (18, 17, 'sp4_r_v_b_24')
// (18, 18, 'neigh_op_tnr_0')
// (18, 18, 'sp4_r_v_b_13')
// (18, 19, 'neigh_op_rgt_0')
// (18, 19, 'sp4_r_v_b_0')
// (18, 20, 'neigh_op_bnr_0')
// (19, 15, 'sp4_h_l_43')
// (19, 15, 'sp4_v_t_37')
// (19, 16, 'sp4_v_b_37')
// (19, 17, 'sp4_v_b_24')
// (19, 18, 'neigh_op_top_0')
// (19, 18, 'sp4_v_b_13')
// (19, 19, 'lutff_0/out')
// (19, 19, 'sp4_v_b_0')
// (19, 20, 'neigh_op_bot_0')
// (20, 18, 'neigh_op_tnl_0')
// (20, 19, 'neigh_op_lft_0')
// (20, 20, 'neigh_op_bnl_0')

reg n970 = 0;
// (15, 15, 'sp4_r_v_b_36')
// (15, 16, 'neigh_op_tnr_6')
// (15, 16, 'sp4_r_v_b_25')
// (15, 17, 'neigh_op_rgt_6')
// (15, 17, 'sp4_r_v_b_12')
// (15, 18, 'neigh_op_bnr_6')
// (15, 18, 'sp4_r_v_b_1')
// (16, 14, 'sp4_h_r_6')
// (16, 14, 'sp4_v_t_36')
// (16, 15, 'sp4_v_b_36')
// (16, 16, 'neigh_op_top_6')
// (16, 16, 'sp4_v_b_25')
// (16, 17, 'lutff_6/out')
// (16, 17, 'sp4_v_b_12')
// (16, 18, 'neigh_op_bot_6')
// (16, 18, 'sp4_v_b_1')
// (17, 14, 'local_g1_3')
// (17, 14, 'lutff_3/in_1')
// (17, 14, 'sp4_h_r_19')
// (17, 16, 'neigh_op_tnl_6')
// (17, 17, 'neigh_op_lft_6')
// (17, 18, 'neigh_op_bnl_6')
// (18, 14, 'sp4_h_r_30')
// (19, 14, 'sp4_h_r_43')
// (20, 14, 'sp4_h_l_43')

reg n971 = 0;
// (15, 15, 'sp4_r_v_b_44')
// (15, 16, 'neigh_op_tnr_2')
// (15, 16, 'sp4_r_v_b_33')
// (15, 17, 'neigh_op_rgt_2')
// (15, 17, 'sp4_r_v_b_20')
// (15, 18, 'neigh_op_bnr_2')
// (15, 18, 'sp4_r_v_b_9')
// (16, 14, 'sp4_v_t_44')
// (16, 15, 'sp4_v_b_44')
// (16, 16, 'neigh_op_top_2')
// (16, 16, 'sp4_v_b_33')
// (16, 17, 'lutff_2/out')
// (16, 17, 'sp4_v_b_20')
// (16, 18, 'neigh_op_bot_2')
// (16, 18, 'sp4_h_r_3')
// (16, 18, 'sp4_v_b_9')
// (17, 16, 'neigh_op_tnl_2')
// (17, 17, 'neigh_op_lft_2')
// (17, 18, 'neigh_op_bnl_2')
// (17, 18, 'sp4_h_r_14')
// (18, 18, 'sp4_h_r_27')
// (19, 18, 'sp4_h_r_38')
// (20, 18, 'sp4_h_l_38')
// (20, 18, 'sp4_h_r_6')
// (21, 18, 'local_g0_3')
// (21, 18, 'lutff_0/in_1')
// (21, 18, 'sp4_h_r_19')
// (22, 18, 'sp4_h_r_30')
// (23, 18, 'sp4_h_r_43')
// (24, 18, 'sp4_h_l_43')

wire n972;
// (15, 16, 'lutff_6/lout')
// (15, 16, 'lutff_7/in_2')

reg n973 = 0;
// (15, 16, 'neigh_op_tnr_0')
// (15, 17, 'neigh_op_rgt_0')
// (15, 18, 'neigh_op_bnr_0')
// (16, 15, 'sp4_r_v_b_41')
// (16, 16, 'neigh_op_top_0')
// (16, 16, 'sp4_r_v_b_28')
// (16, 17, 'lutff_0/out')
// (16, 17, 'sp4_r_v_b_17')
// (16, 18, 'neigh_op_bot_0')
// (16, 18, 'sp4_r_v_b_4')
// (17, 14, 'sp4_v_t_41')
// (17, 15, 'local_g3_1')
// (17, 15, 'lutff_5/in_1')
// (17, 15, 'sp4_v_b_41')
// (17, 16, 'neigh_op_tnl_0')
// (17, 16, 'sp4_v_b_28')
// (17, 17, 'neigh_op_lft_0')
// (17, 17, 'sp4_v_b_17')
// (17, 18, 'neigh_op_bnl_0')
// (17, 18, 'sp4_v_b_4')

reg n974 = 0;
// (15, 16, 'neigh_op_tnr_1')
// (15, 17, 'neigh_op_rgt_1')
// (15, 18, 'neigh_op_bnr_1')
// (16, 15, 'sp4_r_v_b_43')
// (16, 16, 'neigh_op_top_1')
// (16, 16, 'sp4_r_v_b_30')
// (16, 17, 'lutff_1/out')
// (16, 17, 'sp4_r_v_b_19')
// (16, 18, 'neigh_op_bot_1')
// (16, 18, 'sp4_r_v_b_6')
// (17, 14, 'sp4_v_t_43')
// (17, 15, 'local_g3_3')
// (17, 15, 'lutff_7/in_1')
// (17, 15, 'sp4_v_b_43')
// (17, 16, 'neigh_op_tnl_1')
// (17, 16, 'sp4_v_b_30')
// (17, 17, 'neigh_op_lft_1')
// (17, 17, 'sp4_v_b_19')
// (17, 18, 'neigh_op_bnl_1')
// (17, 18, 'sp4_v_b_6')

reg n975 = 0;
// (15, 16, 'neigh_op_tnr_5')
// (15, 17, 'neigh_op_rgt_5')
// (15, 18, 'neigh_op_bnr_5')
// (16, 14, 'sp4_r_v_b_46')
// (16, 15, 'sp4_r_v_b_35')
// (16, 16, 'neigh_op_top_5')
// (16, 16, 'sp4_r_v_b_22')
// (16, 17, 'lutff_5/out')
// (16, 17, 'sp4_r_v_b_11')
// (16, 18, 'neigh_op_bot_5')
// (17, 13, 'sp4_v_t_46')
// (17, 14, 'local_g3_6')
// (17, 14, 'lutff_0/in_1')
// (17, 14, 'sp4_v_b_46')
// (17, 15, 'sp4_v_b_35')
// (17, 16, 'neigh_op_tnl_5')
// (17, 16, 'sp4_v_b_22')
// (17, 17, 'neigh_op_lft_5')
// (17, 17, 'sp4_v_b_11')
// (17, 18, 'neigh_op_bnl_5')

reg n976 = 0;
// (15, 16, 'neigh_op_tnr_7')
// (15, 17, 'neigh_op_rgt_7')
// (15, 18, 'neigh_op_bnr_7')
// (16, 15, 'sp4_r_v_b_39')
// (16, 16, 'neigh_op_top_7')
// (16, 16, 'sp4_r_v_b_26')
// (16, 17, 'lutff_7/out')
// (16, 17, 'sp4_r_v_b_15')
// (16, 18, 'neigh_op_bot_7')
// (16, 18, 'sp4_r_v_b_2')
// (17, 14, 'sp4_v_t_39')
// (17, 15, 'local_g3_7')
// (17, 15, 'lutff_3/in_1')
// (17, 15, 'sp4_v_b_39')
// (17, 16, 'neigh_op_tnl_7')
// (17, 16, 'sp4_v_b_26')
// (17, 17, 'neigh_op_lft_7')
// (17, 17, 'sp4_v_b_15')
// (17, 18, 'neigh_op_bnl_7')
// (17, 18, 'sp4_v_b_2')

reg n977 = 0;
// (15, 16, 'sp4_h_r_4')
// (16, 16, 'sp4_h_r_17')
// (17, 16, 'local_g2_4')
// (17, 16, 'lutff_1/in_3')
// (17, 16, 'sp4_h_r_28')
// (18, 16, 'sp4_h_r_41')
// (19, 16, 'sp4_h_l_41')
// (19, 16, 'sp4_h_r_8')
// (20, 16, 'sp4_h_r_21')
// (21, 16, 'sp4_h_r_32')
// (22, 13, 'sp4_r_v_b_38')
// (22, 14, 'neigh_op_tnr_7')
// (22, 14, 'sp4_r_v_b_27')
// (22, 15, 'neigh_op_rgt_7')
// (22, 15, 'sp4_r_v_b_14')
// (22, 16, 'neigh_op_bnr_7')
// (22, 16, 'sp4_h_r_45')
// (22, 16, 'sp4_r_v_b_3')
// (23, 12, 'sp4_v_t_38')
// (23, 13, 'sp4_v_b_38')
// (23, 14, 'neigh_op_top_7')
// (23, 14, 'sp4_v_b_27')
// (23, 15, 'lutff_7/out')
// (23, 15, 'sp4_v_b_14')
// (23, 16, 'neigh_op_bot_7')
// (23, 16, 'sp4_h_l_45')
// (23, 16, 'sp4_v_b_3')
// (24, 14, 'neigh_op_tnl_7')
// (24, 15, 'neigh_op_lft_7')
// (24, 16, 'neigh_op_bnl_7')

reg n978 = 0;
// (15, 16, 'sp4_h_r_9')
// (16, 16, 'sp4_h_r_20')
// (17, 16, 'local_g3_1')
// (17, 16, 'lutff_1/in_1')
// (17, 16, 'sp4_h_r_33')
// (18, 16, 'sp4_h_r_44')
// (19, 16, 'sp4_h_l_44')
// (19, 16, 'sp4_h_r_6')
// (20, 16, 'sp4_h_r_19')
// (21, 16, 'sp4_h_r_30')
// (22, 13, 'neigh_op_tnr_7')
// (22, 13, 'sp4_r_v_b_43')
// (22, 14, 'neigh_op_rgt_7')
// (22, 14, 'sp4_r_v_b_30')
// (22, 15, 'neigh_op_bnr_7')
// (22, 15, 'sp4_r_v_b_19')
// (22, 16, 'sp4_h_r_43')
// (22, 16, 'sp4_r_v_b_6')
// (23, 12, 'sp4_v_t_43')
// (23, 13, 'neigh_op_top_7')
// (23, 13, 'sp4_v_b_43')
// (23, 14, 'lutff_7/out')
// (23, 14, 'sp4_v_b_30')
// (23, 15, 'neigh_op_bot_7')
// (23, 15, 'sp4_v_b_19')
// (23, 16, 'sp4_h_l_43')
// (23, 16, 'sp4_v_b_6')
// (24, 13, 'neigh_op_tnl_7')
// (24, 14, 'neigh_op_lft_7')
// (24, 15, 'neigh_op_bnl_7')

reg n979 = 0;
// (15, 17, 'neigh_op_tnr_0')
// (15, 18, 'neigh_op_rgt_0')
// (15, 19, 'neigh_op_bnr_0')
// (16, 16, 'sp4_r_v_b_41')
// (16, 17, 'neigh_op_top_0')
// (16, 17, 'sp4_r_v_b_28')
// (16, 18, 'lutff_0/out')
// (16, 18, 'sp4_r_v_b_17')
// (16, 19, 'neigh_op_bot_0')
// (16, 19, 'sp4_r_v_b_4')
// (16, 20, 'sp4_r_v_b_42')
// (16, 21, 'sp4_r_v_b_31')
// (16, 22, 'sp4_r_v_b_18')
// (16, 23, 'sp4_r_v_b_7')
// (17, 15, 'sp4_v_t_41')
// (17, 16, 'sp4_v_b_41')
// (17, 17, 'neigh_op_tnl_0')
// (17, 17, 'sp4_v_b_28')
// (17, 18, 'local_g1_1')
// (17, 18, 'lutff_0/in_2')
// (17, 18, 'neigh_op_lft_0')
// (17, 18, 'sp4_v_b_17')
// (17, 19, 'neigh_op_bnl_0')
// (17, 19, 'sp4_v_b_4')
// (17, 19, 'sp4_v_t_42')
// (17, 20, 'sp4_v_b_42')
// (17, 21, 'sp4_v_b_31')
// (17, 22, 'local_g1_2')
// (17, 22, 'lutff_0/in_3')
// (17, 22, 'sp4_v_b_18')
// (17, 23, 'sp4_v_b_7')

reg n980 = 0;
// (15, 17, 'neigh_op_tnr_2')
// (15, 18, 'neigh_op_rgt_2')
// (15, 18, 'sp4_h_r_9')
// (15, 19, 'neigh_op_bnr_2')
// (15, 22, 'sp4_h_r_2')
// (16, 17, 'neigh_op_top_2')
// (16, 18, 'lutff_2/out')
// (16, 18, 'sp4_h_r_20')
// (16, 19, 'neigh_op_bot_2')
// (16, 22, 'sp4_h_r_15')
// (17, 17, 'neigh_op_tnl_2')
// (17, 18, 'local_g3_1')
// (17, 18, 'lutff_2/in_2')
// (17, 18, 'neigh_op_lft_2')
// (17, 18, 'sp4_h_r_33')
// (17, 19, 'neigh_op_bnl_2')
// (17, 22, 'local_g3_2')
// (17, 22, 'lutff_2/in_3')
// (17, 22, 'sp4_h_r_26')
// (18, 18, 'sp4_h_r_44')
// (18, 19, 'sp4_r_v_b_39')
// (18, 20, 'sp4_r_v_b_26')
// (18, 21, 'sp4_r_v_b_15')
// (18, 22, 'sp4_h_r_39')
// (18, 22, 'sp4_r_v_b_2')
// (19, 18, 'sp4_h_l_44')
// (19, 18, 'sp4_v_t_39')
// (19, 19, 'sp4_v_b_39')
// (19, 20, 'sp4_v_b_26')
// (19, 21, 'sp4_v_b_15')
// (19, 22, 'sp4_h_l_39')
// (19, 22, 'sp4_v_b_2')

reg n981 = 0;
// (15, 17, 'neigh_op_tnr_3')
// (15, 18, 'neigh_op_rgt_3')
// (15, 19, 'neigh_op_bnr_3')
// (16, 17, 'neigh_op_top_3')
// (16, 18, 'lutff_3/out')
// (16, 18, 'sp4_r_v_b_39')
// (16, 19, 'neigh_op_bot_3')
// (16, 19, 'sp4_r_v_b_26')
// (16, 20, 'sp4_r_v_b_15')
// (16, 21, 'sp4_r_v_b_2')
// (16, 22, 'sp4_r_v_b_40')
// (16, 23, 'sp4_r_v_b_29')
// (16, 24, 'sp4_r_v_b_16')
// (16, 25, 'sp4_r_v_b_5')
// (17, 17, 'neigh_op_tnl_3')
// (17, 17, 'sp4_v_t_39')
// (17, 18, 'local_g0_3')
// (17, 18, 'lutff_3/in_2')
// (17, 18, 'neigh_op_lft_3')
// (17, 18, 'sp4_v_b_39')
// (17, 19, 'neigh_op_bnl_3')
// (17, 19, 'sp4_v_b_26')
// (17, 20, 'sp4_v_b_15')
// (17, 21, 'sp4_v_b_2')
// (17, 21, 'sp4_v_t_40')
// (17, 22, 'local_g2_0')
// (17, 22, 'lutff_3/in_3')
// (17, 22, 'sp4_v_b_40')
// (17, 23, 'sp4_v_b_29')
// (17, 24, 'sp4_v_b_16')
// (17, 25, 'sp4_v_b_5')

reg n982 = 0;
// (15, 17, 'neigh_op_tnr_4')
// (15, 18, 'neigh_op_rgt_4')
// (15, 19, 'neigh_op_bnr_4')
// (16, 17, 'neigh_op_top_4')
// (16, 17, 'sp4_r_v_b_36')
// (16, 18, 'lutff_4/out')
// (16, 18, 'sp4_h_r_8')
// (16, 18, 'sp4_r_v_b_25')
// (16, 19, 'neigh_op_bot_4')
// (16, 19, 'sp4_r_v_b_12')
// (16, 20, 'sp4_r_v_b_1')
// (16, 21, 'sp4_r_v_b_41')
// (16, 22, 'sp4_r_v_b_28')
// (16, 23, 'sp4_r_v_b_17')
// (16, 24, 'sp4_r_v_b_4')
// (17, 16, 'sp4_v_t_36')
// (17, 17, 'neigh_op_tnl_4')
// (17, 17, 'sp4_v_b_36')
// (17, 18, 'local_g0_5')
// (17, 18, 'lutff_4/in_1')
// (17, 18, 'neigh_op_lft_4')
// (17, 18, 'sp4_h_r_21')
// (17, 18, 'sp4_v_b_25')
// (17, 19, 'neigh_op_bnl_4')
// (17, 19, 'sp4_v_b_12')
// (17, 20, 'sp4_v_b_1')
// (17, 20, 'sp4_v_t_41')
// (17, 21, 'sp4_v_b_41')
// (17, 22, 'local_g3_4')
// (17, 22, 'lutff_4/in_3')
// (17, 22, 'sp4_v_b_28')
// (17, 23, 'sp4_v_b_17')
// (17, 24, 'sp4_v_b_4')
// (18, 18, 'sp4_h_r_32')
// (19, 18, 'sp4_h_r_45')
// (20, 18, 'sp4_h_l_45')

reg n983 = 0;
// (15, 17, 'neigh_op_tnr_7')
// (15, 18, 'neigh_op_rgt_7')
// (15, 19, 'neigh_op_bnr_7')
// (16, 17, 'neigh_op_top_7')
// (16, 18, 'lutff_7/out')
// (16, 18, 'sp4_r_v_b_47')
// (16, 19, 'neigh_op_bot_7')
// (16, 19, 'sp4_r_v_b_34')
// (16, 20, 'sp4_r_v_b_23')
// (16, 21, 'sp4_r_v_b_10')
// (16, 22, 'sp4_r_v_b_36')
// (16, 23, 'sp4_r_v_b_25')
// (16, 24, 'sp4_r_v_b_12')
// (16, 25, 'sp4_r_v_b_1')
// (17, 17, 'neigh_op_tnl_7')
// (17, 17, 'sp4_v_t_47')
// (17, 18, 'local_g1_7')
// (17, 18, 'lutff_7/in_1')
// (17, 18, 'neigh_op_lft_7')
// (17, 18, 'sp4_v_b_47')
// (17, 19, 'neigh_op_bnl_7')
// (17, 19, 'sp4_v_b_34')
// (17, 20, 'sp4_v_b_23')
// (17, 21, 'sp4_v_b_10')
// (17, 21, 'sp4_v_t_36')
// (17, 22, 'local_g2_4')
// (17, 22, 'lutff_7/in_3')
// (17, 22, 'sp4_v_b_36')
// (17, 23, 'sp4_v_b_25')
// (17, 24, 'sp4_v_b_12')
// (17, 25, 'sp4_v_b_1')

reg n984 = 0;
// (15, 17, 'sp4_h_r_0')
// (16, 17, 'sp4_h_r_13')
// (17, 17, 'local_g2_0')
// (17, 17, 'lutff_5/in_3')
// (17, 17, 'sp4_h_r_24')
// (18, 17, 'sp4_h_r_37')
// (19, 17, 'sp4_h_l_37')
// (19, 17, 'sp4_h_r_9')
// (20, 17, 'sp4_h_r_20')
// (21, 17, 'sp4_h_r_33')
// (22, 17, 'sp4_h_r_44')
// (23, 17, 'sp4_h_l_44')
// (23, 17, 'sp4_h_r_1')
// (24, 17, 'sp4_h_r_12')
// (25, 16, 'neigh_op_tnr_2')
// (25, 17, 'neigh_op_rgt_2')
// (25, 17, 'sp4_h_r_25')
// (25, 18, 'neigh_op_bnr_2')
// (26, 16, 'neigh_op_top_2')
// (26, 17, 'lutff_2/out')
// (26, 17, 'sp4_h_r_36')
// (26, 18, 'neigh_op_bot_2')
// (27, 16, 'neigh_op_tnl_2')
// (27, 17, 'neigh_op_lft_2')
// (27, 17, 'sp4_h_l_36')
// (27, 18, 'neigh_op_bnl_2')

wire n985;
// (15, 17, 'sp4_h_r_3')
// (16, 17, 'sp4_h_r_14')
// (17, 17, 'local_g3_3')
// (17, 17, 'lutff_global/cen')
// (17, 17, 'sp4_h_r_27')
// (18, 17, 'sp4_h_r_38')
// (18, 18, 'sp4_r_v_b_38')
// (18, 19, 'neigh_op_tnr_7')
// (18, 19, 'sp4_r_v_b_27')
// (18, 19, 'sp4_r_v_b_43')
// (18, 20, 'neigh_op_rgt_7')
// (18, 20, 'sp4_r_v_b_14')
// (18, 20, 'sp4_r_v_b_30')
// (18, 21, 'neigh_op_bnr_7')
// (18, 21, 'sp4_r_v_b_19')
// (18, 21, 'sp4_r_v_b_3')
// (18, 22, 'sp4_r_v_b_6')
// (19, 17, 'sp4_h_l_38')
// (19, 17, 'sp4_v_t_38')
// (19, 18, 'sp4_v_b_38')
// (19, 18, 'sp4_v_t_43')
// (19, 19, 'local_g3_3')
// (19, 19, 'lutff_global/cen')
// (19, 19, 'neigh_op_top_7')
// (19, 19, 'sp4_v_b_27')
// (19, 19, 'sp4_v_b_43')
// (19, 20, 'lutff_7/out')
// (19, 20, 'sp4_v_b_14')
// (19, 20, 'sp4_v_b_30')
// (19, 21, 'neigh_op_bot_7')
// (19, 21, 'sp4_v_b_19')
// (19, 21, 'sp4_v_b_3')
// (19, 22, 'sp4_v_b_6')
// (20, 19, 'neigh_op_tnl_7')
// (20, 20, 'neigh_op_lft_7')
// (20, 21, 'neigh_op_bnl_7')

reg n986 = 0;
// (15, 17, 'sp4_h_r_9')
// (16, 17, 'sp4_h_r_20')
// (17, 17, 'local_g3_1')
// (17, 17, 'lutff_3/in_3')
// (17, 17, 'sp4_h_r_33')
// (18, 10, 'neigh_op_tnr_0')
// (18, 10, 'sp4_r_v_b_45')
// (18, 11, 'neigh_op_rgt_0')
// (18, 11, 'sp4_r_v_b_32')
// (18, 12, 'neigh_op_bnr_0')
// (18, 12, 'sp4_r_v_b_21')
// (18, 13, 'sp4_r_v_b_8')
// (18, 14, 'sp4_r_v_b_41')
// (18, 15, 'sp4_r_v_b_28')
// (18, 16, 'sp4_r_v_b_17')
// (18, 17, 'sp4_h_r_44')
// (18, 17, 'sp4_r_v_b_4')
// (19, 9, 'sp4_v_t_45')
// (19, 10, 'neigh_op_top_0')
// (19, 10, 'sp4_v_b_45')
// (19, 11, 'lutff_0/out')
// (19, 11, 'sp4_v_b_32')
// (19, 12, 'neigh_op_bot_0')
// (19, 12, 'sp4_v_b_21')
// (19, 13, 'sp4_v_b_8')
// (19, 13, 'sp4_v_t_41')
// (19, 14, 'sp4_v_b_41')
// (19, 15, 'sp4_v_b_28')
// (19, 16, 'sp4_v_b_17')
// (19, 17, 'sp4_h_l_44')
// (19, 17, 'sp4_v_b_4')
// (20, 10, 'neigh_op_tnl_0')
// (20, 11, 'neigh_op_lft_0')
// (20, 12, 'neigh_op_bnl_0')

reg n987 = 0;
// (15, 18, 'neigh_op_tnr_1')
// (15, 19, 'neigh_op_rgt_1')
// (15, 20, 'neigh_op_bnr_1')
// (16, 17, 'sp4_r_v_b_43')
// (16, 18, 'neigh_op_top_1')
// (16, 18, 'sp4_r_v_b_30')
// (16, 19, 'lutff_1/out')
// (16, 19, 'sp4_r_v_b_19')
// (16, 20, 'neigh_op_bot_1')
// (16, 20, 'sp4_r_v_b_6')
// (16, 21, 'sp4_r_v_b_39')
// (16, 22, 'sp4_r_v_b_26')
// (16, 23, 'sp4_r_v_b_15')
// (16, 24, 'sp4_r_v_b_2')
// (17, 16, 'sp4_v_t_43')
// (17, 17, 'sp4_v_b_43')
// (17, 18, 'neigh_op_tnl_1')
// (17, 18, 'sp4_v_b_30')
// (17, 19, 'local_g0_1')
// (17, 19, 'lutff_3/in_2')
// (17, 19, 'neigh_op_lft_1')
// (17, 19, 'sp4_v_b_19')
// (17, 20, 'neigh_op_bnl_1')
// (17, 20, 'sp4_v_b_6')
// (17, 20, 'sp4_v_t_39')
// (17, 21, 'sp4_v_b_39')
// (17, 22, 'sp4_v_b_26')
// (17, 23, 'local_g1_7')
// (17, 23, 'lutff_3/in_3')
// (17, 23, 'sp4_v_b_15')
// (17, 24, 'sp4_v_b_2')

reg n988 = 0;
// (15, 18, 'neigh_op_tnr_3')
// (15, 19, 'neigh_op_rgt_3')
// (15, 20, 'neigh_op_bnr_3')
// (16, 17, 'sp4_r_v_b_47')
// (16, 18, 'neigh_op_top_3')
// (16, 18, 'sp4_r_v_b_34')
// (16, 19, 'lutff_3/out')
// (16, 19, 'sp4_r_v_b_23')
// (16, 20, 'neigh_op_bot_3')
// (16, 20, 'sp4_r_v_b_10')
// (16, 21, 'sp4_r_v_b_43')
// (16, 22, 'sp4_r_v_b_30')
// (16, 23, 'sp4_r_v_b_19')
// (16, 24, 'sp4_r_v_b_6')
// (17, 16, 'sp4_v_t_47')
// (17, 17, 'sp4_v_b_47')
// (17, 18, 'neigh_op_tnl_3')
// (17, 18, 'sp4_v_b_34')
// (17, 19, 'local_g1_3')
// (17, 19, 'lutff_5/in_1')
// (17, 19, 'neigh_op_lft_3')
// (17, 19, 'sp4_v_b_23')
// (17, 20, 'neigh_op_bnl_3')
// (17, 20, 'sp4_v_b_10')
// (17, 20, 'sp4_v_t_43')
// (17, 21, 'sp4_v_b_43')
// (17, 22, 'sp4_v_b_30')
// (17, 23, 'local_g1_3')
// (17, 23, 'lutff_5/in_3')
// (17, 23, 'sp4_v_b_19')
// (17, 24, 'sp4_v_b_6')

reg n989 = 0;
// (15, 18, 'neigh_op_tnr_4')
// (15, 19, 'neigh_op_rgt_4')
// (15, 20, 'neigh_op_bnr_4')
// (16, 18, 'neigh_op_top_4')
// (16, 19, 'lutff_4/out')
// (16, 19, 'sp4_h_r_8')
// (16, 19, 'sp4_r_v_b_41')
// (16, 20, 'neigh_op_bot_4')
// (16, 20, 'sp4_r_v_b_28')
// (16, 21, 'sp4_r_v_b_17')
// (16, 22, 'sp4_r_v_b_4')
// (16, 23, 'sp4_r_v_b_42')
// (16, 24, 'sp4_r_v_b_31')
// (16, 25, 'sp4_r_v_b_18')
// (16, 26, 'sp4_r_v_b_7')
// (17, 18, 'neigh_op_tnl_4')
// (17, 18, 'sp4_v_t_41')
// (17, 19, 'local_g0_5')
// (17, 19, 'lutff_6/in_1')
// (17, 19, 'neigh_op_lft_4')
// (17, 19, 'sp4_h_r_21')
// (17, 19, 'sp4_v_b_41')
// (17, 20, 'neigh_op_bnl_4')
// (17, 20, 'sp4_v_b_28')
// (17, 21, 'sp4_v_b_17')
// (17, 22, 'sp4_v_b_4')
// (17, 22, 'sp4_v_t_42')
// (17, 23, 'local_g3_2')
// (17, 23, 'lutff_6/in_3')
// (17, 23, 'sp4_v_b_42')
// (17, 24, 'sp4_v_b_31')
// (17, 25, 'sp4_v_b_18')
// (17, 26, 'sp4_v_b_7')
// (18, 19, 'sp4_h_r_32')
// (19, 19, 'sp4_h_r_45')
// (20, 19, 'sp4_h_l_45')

reg n990 = 0;
// (15, 18, 'neigh_op_tnr_5')
// (15, 19, 'neigh_op_rgt_5')
// (15, 20, 'neigh_op_bnr_5')
// (16, 18, 'neigh_op_top_5')
// (16, 19, 'lutff_5/out')
// (16, 19, 'sp4_r_v_b_43')
// (16, 20, 'neigh_op_bot_5')
// (16, 20, 'sp4_r_v_b_30')
// (16, 21, 'sp4_r_v_b_19')
// (16, 22, 'sp4_r_v_b_6')
// (16, 23, 'sp4_r_v_b_44')
// (16, 24, 'sp4_r_v_b_33')
// (16, 25, 'sp4_r_v_b_20')
// (16, 26, 'sp4_r_v_b_9')
// (17, 18, 'neigh_op_tnl_5')
// (17, 18, 'sp4_v_t_43')
// (17, 19, 'local_g1_5')
// (17, 19, 'lutff_7/in_1')
// (17, 19, 'neigh_op_lft_5')
// (17, 19, 'sp4_v_b_43')
// (17, 20, 'neigh_op_bnl_5')
// (17, 20, 'sp4_v_b_30')
// (17, 21, 'sp4_v_b_19')
// (17, 22, 'sp4_v_b_6')
// (17, 22, 'sp4_v_t_44')
// (17, 23, 'local_g2_4')
// (17, 23, 'lutff_7/in_3')
// (17, 23, 'sp4_v_b_44')
// (17, 24, 'sp4_v_b_33')
// (17, 25, 'sp4_v_b_20')
// (17, 26, 'sp4_v_b_9')

reg n991 = 0;
// (15, 18, 'neigh_op_tnr_6')
// (15, 19, 'neigh_op_rgt_6')
// (15, 19, 'sp4_h_r_1')
// (15, 20, 'neigh_op_bnr_6')
// (15, 23, 'sp4_h_r_11')
// (16, 18, 'neigh_op_top_6')
// (16, 19, 'lutff_6/out')
// (16, 19, 'sp4_h_r_12')
// (16, 20, 'neigh_op_bot_6')
// (16, 23, 'sp4_h_r_22')
// (17, 18, 'neigh_op_tnl_6')
// (17, 19, 'local_g3_1')
// (17, 19, 'lutff_0/in_2')
// (17, 19, 'neigh_op_lft_6')
// (17, 19, 'sp4_h_r_25')
// (17, 20, 'neigh_op_bnl_6')
// (17, 23, 'local_g2_3')
// (17, 23, 'lutff_0/in_3')
// (17, 23, 'sp4_h_r_35')
// (18, 19, 'sp4_h_r_36')
// (18, 20, 'sp4_r_v_b_43')
// (18, 21, 'sp4_r_v_b_30')
// (18, 22, 'sp4_r_v_b_19')
// (18, 23, 'sp4_h_r_46')
// (18, 23, 'sp4_r_v_b_6')
// (19, 19, 'sp4_h_l_36')
// (19, 19, 'sp4_v_t_43')
// (19, 20, 'sp4_v_b_43')
// (19, 21, 'sp4_v_b_30')
// (19, 22, 'sp4_v_b_19')
// (19, 23, 'sp4_h_l_46')
// (19, 23, 'sp4_v_b_6')

reg n992 = 0;
// (15, 18, 'neigh_op_tnr_7')
// (15, 19, 'neigh_op_rgt_7')
// (15, 20, 'neigh_op_bnr_7')
// (16, 18, 'neigh_op_top_7')
// (16, 18, 'sp4_r_v_b_42')
// (16, 19, 'lutff_7/out')
// (16, 19, 'sp4_r_v_b_31')
// (16, 20, 'neigh_op_bot_7')
// (16, 20, 'sp4_r_v_b_18')
// (16, 21, 'sp4_r_v_b_7')
// (16, 22, 'sp4_r_v_b_47')
// (16, 23, 'sp4_r_v_b_34')
// (16, 24, 'sp4_r_v_b_23')
// (16, 25, 'sp4_r_v_b_10')
// (17, 17, 'sp4_v_t_42')
// (17, 18, 'neigh_op_tnl_7')
// (17, 18, 'sp4_v_b_42')
// (17, 19, 'local_g0_7')
// (17, 19, 'lutff_1/in_2')
// (17, 19, 'neigh_op_lft_7')
// (17, 19, 'sp4_v_b_31')
// (17, 20, 'neigh_op_bnl_7')
// (17, 20, 'sp4_v_b_18')
// (17, 21, 'sp4_v_b_7')
// (17, 21, 'sp4_v_t_47')
// (17, 22, 'sp4_v_b_47')
// (17, 23, 'local_g2_2')
// (17, 23, 'lutff_1/in_3')
// (17, 23, 'sp4_v_b_34')
// (17, 24, 'sp4_v_b_23')
// (17, 25, 'sp4_v_b_10')

wire n993;
// (15, 18, 'sp4_r_v_b_36')
// (15, 19, 'sp4_r_v_b_25')
// (15, 20, 'sp4_r_v_b_12')
// (15, 21, 'sp4_r_v_b_1')
// (16, 17, 'sp4_h_r_1')
// (16, 17, 'sp4_v_t_36')
// (16, 18, 'sp4_v_b_36')
// (16, 19, 'sp4_v_b_25')
// (16, 20, 'neigh_op_tnr_6')
// (16, 20, 'sp4_v_b_12')
// (16, 21, 'neigh_op_rgt_6')
// (16, 21, 'sp4_h_r_1')
// (16, 21, 'sp4_v_b_1')
// (16, 22, 'neigh_op_bnr_6')
// (17, 17, 'sp4_h_r_12')
// (17, 20, 'neigh_op_top_6')
// (17, 21, 'lutff_6/out')
// (17, 21, 'sp4_h_r_12')
// (17, 22, 'neigh_op_bot_6')
// (18, 17, 'sp4_h_r_25')
// (18, 20, 'neigh_op_tnl_6')
// (18, 21, 'neigh_op_lft_6')
// (18, 21, 'sp4_h_r_25')
// (18, 22, 'neigh_op_bnl_6')
// (19, 17, 'local_g3_4')
// (19, 17, 'lutff_4/in_1')
// (19, 17, 'sp4_h_r_36')
// (19, 21, 'sp4_h_r_36')
// (20, 17, 'sp4_h_l_36')
// (20, 21, 'sp4_h_l_36')

reg n994 = 0;
// (15, 19, 'neigh_op_tnr_0')
// (15, 19, 'sp4_r_v_b_45')
// (15, 20, 'neigh_op_rgt_0')
// (15, 20, 'sp4_r_v_b_32')
// (15, 21, 'neigh_op_bnr_0')
// (15, 21, 'sp4_r_v_b_21')
// (15, 22, 'sp4_r_v_b_8')
// (16, 18, 'sp4_v_t_45')
// (16, 19, 'neigh_op_top_0')
// (16, 19, 'sp4_v_b_45')
// (16, 20, 'local_g0_0')
// (16, 20, 'lutff_0/in_0')
// (16, 20, 'lutff_0/out')
// (16, 20, 'sp4_v_b_32')
// (16, 21, 'neigh_op_bot_0')
// (16, 21, 'sp4_v_b_21')
// (16, 22, 'sp4_h_r_2')
// (16, 22, 'sp4_v_b_8')
// (17, 19, 'neigh_op_tnl_0')
// (17, 20, 'neigh_op_lft_0')
// (17, 21, 'neigh_op_bnl_0')
// (17, 22, 'sp4_h_r_15')
// (18, 22, 'sp4_h_r_26')
// (19, 22, 'sp4_h_r_39')
// (20, 22, 'local_g0_2')
// (20, 22, 'lutff_7/in_1')
// (20, 22, 'sp4_h_l_39')
// (20, 22, 'sp4_h_r_2')
// (21, 22, 'sp4_h_r_15')
// (22, 22, 'sp4_h_r_26')
// (23, 22, 'sp4_h_r_39')
// (24, 22, 'sp4_h_l_39')

wire n995;
// (15, 19, 'neigh_op_tnr_4')
// (15, 20, 'neigh_op_rgt_4')
// (15, 20, 'sp4_r_v_b_40')
// (15, 20, 'sp4_r_v_b_46')
// (15, 21, 'neigh_op_bnr_4')
// (15, 21, 'sp4_r_v_b_29')
// (15, 21, 'sp4_r_v_b_35')
// (15, 22, 'sp4_r_v_b_16')
// (15, 22, 'sp4_r_v_b_22')
// (15, 23, 'sp4_r_v_b_11')
// (15, 23, 'sp4_r_v_b_5')
// (16, 19, 'neigh_op_top_4')
// (16, 19, 'sp4_h_r_5')
// (16, 19, 'sp4_v_t_40')
// (16, 19, 'sp4_v_t_46')
// (16, 20, 'lutff_4/out')
// (16, 20, 'sp4_v_b_40')
// (16, 20, 'sp4_v_b_46')
// (16, 21, 'local_g3_3')
// (16, 21, 'lutff_global/cen')
// (16, 21, 'neigh_op_bot_4')
// (16, 21, 'sp4_v_b_29')
// (16, 21, 'sp4_v_b_35')
// (16, 22, 'sp4_v_b_16')
// (16, 22, 'sp4_v_b_22')
// (16, 23, 'sp4_v_b_11')
// (16, 23, 'sp4_v_b_5')
// (17, 19, 'neigh_op_tnl_4')
// (17, 19, 'sp4_h_r_16')
// (17, 20, 'neigh_op_lft_4')
// (17, 21, 'neigh_op_bnl_4')
// (18, 19, 'sp4_h_r_29')
// (19, 19, 'sp4_h_r_40')
// (20, 19, 'sp4_h_l_40')

wire n996;
// (15, 19, 'neigh_op_tnr_7')
// (15, 20, 'neigh_op_rgt_7')
// (15, 20, 'sp4_h_r_3')
// (15, 21, 'neigh_op_bnr_7')
// (16, 19, 'neigh_op_top_7')
// (16, 20, 'lutff_7/out')
// (16, 20, 'sp4_h_r_14')
// (16, 21, 'neigh_op_bot_7')
// (17, 19, 'neigh_op_tnl_7')
// (17, 20, 'neigh_op_lft_7')
// (17, 20, 'sp4_h_r_27')
// (17, 21, 'neigh_op_bnl_7')
// (18, 20, 'sp4_h_r_38')
// (19, 20, 'sp4_h_l_38')
// (19, 20, 'sp4_h_r_6')
// (20, 20, 'local_g1_3')
// (20, 20, 'lutff_global/cen')
// (20, 20, 'sp4_h_r_19')
// (21, 20, 'sp4_h_r_30')
// (22, 20, 'sp4_h_r_43')
// (23, 20, 'sp4_h_l_43')

wire n997;
// (15, 20, 'lutff_7/cout')
// (15, 21, 'carry_in')
// (15, 21, 'carry_in_mux')

reg n998 = 0;
// (15, 20, 'neigh_op_tnr_0')
// (15, 21, 'local_g2_0')
// (15, 21, 'lutff_2/in_0')
// (15, 21, 'neigh_op_rgt_0')
// (15, 22, 'neigh_op_bnr_0')
// (16, 20, 'neigh_op_top_0')
// (16, 21, 'lutff_0/out')
// (16, 22, 'neigh_op_bot_0')
// (17, 20, 'neigh_op_tnl_0')
// (17, 21, 'neigh_op_lft_0')
// (17, 22, 'neigh_op_bnl_0')

reg n999 = 0;
// (15, 20, 'neigh_op_tnr_1')
// (15, 21, 'local_g2_1')
// (15, 21, 'lutff_3/in_0')
// (15, 21, 'neigh_op_rgt_1')
// (15, 22, 'neigh_op_bnr_1')
// (16, 20, 'neigh_op_top_1')
// (16, 21, 'lutff_1/out')
// (16, 22, 'neigh_op_bot_1')
// (17, 20, 'neigh_op_tnl_1')
// (17, 21, 'neigh_op_lft_1')
// (17, 22, 'neigh_op_bnl_1')

reg n1000 = 0;
// (15, 20, 'neigh_op_tnr_2')
// (15, 21, 'local_g3_2')
// (15, 21, 'lutff_4/in_3')
// (15, 21, 'neigh_op_rgt_2')
// (15, 22, 'neigh_op_bnr_2')
// (16, 20, 'neigh_op_top_2')
// (16, 21, 'lutff_2/out')
// (16, 22, 'neigh_op_bot_2')
// (17, 20, 'neigh_op_tnl_2')
// (17, 21, 'neigh_op_lft_2')
// (17, 22, 'neigh_op_bnl_2')

reg n1001 = 0;
// (15, 20, 'neigh_op_tnr_3')
// (15, 21, 'local_g3_3')
// (15, 21, 'lutff_5/in_3')
// (15, 21, 'neigh_op_rgt_3')
// (15, 22, 'neigh_op_bnr_3')
// (16, 20, 'neigh_op_top_3')
// (16, 21, 'lutff_3/out')
// (16, 22, 'neigh_op_bot_3')
// (17, 20, 'neigh_op_tnl_3')
// (17, 21, 'neigh_op_lft_3')
// (17, 22, 'neigh_op_bnl_3')

reg n1002 = 0;
// (15, 20, 'neigh_op_tnr_4')
// (15, 21, 'local_g2_4')
// (15, 21, 'lutff_6/in_0')
// (15, 21, 'neigh_op_rgt_4')
// (15, 22, 'neigh_op_bnr_4')
// (16, 20, 'neigh_op_top_4')
// (16, 21, 'lutff_4/out')
// (16, 22, 'neigh_op_bot_4')
// (17, 20, 'neigh_op_tnl_4')
// (17, 21, 'neigh_op_lft_4')
// (17, 22, 'neigh_op_bnl_4')

reg n1003 = 0;
// (15, 20, 'neigh_op_tnr_5')
// (15, 21, 'local_g2_5')
// (15, 21, 'lutff_7/in_0')
// (15, 21, 'neigh_op_rgt_5')
// (15, 22, 'neigh_op_bnr_5')
// (16, 20, 'neigh_op_top_5')
// (16, 21, 'lutff_5/out')
// (16, 22, 'neigh_op_bot_5')
// (17, 20, 'neigh_op_tnl_5')
// (17, 21, 'neigh_op_lft_5')
// (17, 22, 'neigh_op_bnl_5')

reg n1004 = 0;
// (15, 20, 'neigh_op_tnr_6')
// (15, 21, 'local_g3_6')
// (15, 21, 'lutff_0/in_3')
// (15, 21, 'neigh_op_rgt_6')
// (15, 22, 'neigh_op_bnr_6')
// (16, 20, 'neigh_op_top_6')
// (16, 21, 'lutff_6/out')
// (16, 22, 'neigh_op_bot_6')
// (17, 20, 'neigh_op_tnl_6')
// (17, 21, 'neigh_op_lft_6')
// (17, 22, 'neigh_op_bnl_6')

reg n1005 = 0;
// (15, 20, 'neigh_op_tnr_7')
// (15, 21, 'local_g3_7')
// (15, 21, 'lutff_1/in_3')
// (15, 21, 'neigh_op_rgt_7')
// (15, 22, 'neigh_op_bnr_7')
// (16, 20, 'neigh_op_top_7')
// (16, 21, 'lutff_7/out')
// (16, 22, 'neigh_op_bot_7')
// (17, 20, 'neigh_op_tnl_7')
// (17, 21, 'neigh_op_lft_7')
// (17, 22, 'neigh_op_bnl_7')

wire n1006;
// (15, 21, 'lutff_7/cout')
// (15, 22, 'carry_in')
// (15, 22, 'carry_in_mux')

reg io_33_30_0 = 0;
// (15, 21, 'neigh_op_tnr_0')
// (15, 22, 'neigh_op_rgt_0')
// (15, 23, 'neigh_op_bnr_0')
// (16, 18, 'sp12_v_t_23')
// (16, 19, 'sp12_v_b_23')
// (16, 20, 'sp12_v_b_20')
// (16, 21, 'neigh_op_top_0')
// (16, 21, 'sp12_v_b_19')
// (16, 22, 'lutff_0/out')
// (16, 22, 'sp12_v_b_16')
// (16, 23, 'neigh_op_bot_0')
// (16, 23, 'sp12_v_b_15')
// (16, 24, 'sp12_v_b_12')
// (16, 25, 'sp12_v_b_11')
// (16, 26, 'sp12_v_b_8')
// (16, 27, 'sp12_v_b_7')
// (16, 28, 'sp12_v_b_4')
// (16, 29, 'sp12_v_b_3')
// (16, 30, 'sp12_h_r_0')
// (16, 30, 'sp12_v_b_0')
// (17, 21, 'neigh_op_tnl_0')
// (17, 22, 'neigh_op_lft_0')
// (17, 23, 'neigh_op_bnl_0')
// (17, 30, 'sp12_h_r_3')
// (18, 30, 'sp12_h_r_4')
// (19, 30, 'sp12_h_r_7')
// (20, 30, 'sp12_h_r_8')
// (21, 30, 'sp12_h_r_11')
// (22, 30, 'sp12_h_r_12')
// (23, 30, 'sp12_h_r_15')
// (24, 30, 'sp12_h_r_16')
// (25, 30, 'sp12_h_r_19')
// (26, 30, 'sp12_h_r_20')
// (27, 30, 'sp12_h_r_23')
// (28, 30, 'sp12_h_l_23')
// (28, 30, 'sp12_h_r_0')
// (29, 30, 'sp12_h_r_3')
// (30, 30, 'sp12_h_r_4')
// (31, 30, 'sp12_h_r_7')
// (32, 30, 'sp12_h_r_8')
// (33, 30, 'io_0/D_OUT_0')
// (33, 30, 'io_0/PAD')
// (33, 30, 'local_g0_0')
// (33, 30, 'span12_horz_8')

reg io_33_30_1 = 0;
// (15, 21, 'neigh_op_tnr_1')
// (15, 22, 'neigh_op_rgt_1')
// (15, 23, 'neigh_op_bnr_1')
// (16, 19, 'sp12_v_t_22')
// (16, 20, 'sp12_v_b_22')
// (16, 21, 'neigh_op_top_1')
// (16, 21, 'sp12_v_b_21')
// (16, 22, 'lutff_1/out')
// (16, 22, 'sp12_v_b_18')
// (16, 23, 'neigh_op_bot_1')
// (16, 23, 'sp12_v_b_17')
// (16, 24, 'sp12_v_b_14')
// (16, 25, 'sp12_v_b_13')
// (16, 26, 'sp12_v_b_10')
// (16, 27, 'sp12_v_b_9')
// (16, 28, 'sp12_v_b_6')
// (16, 29, 'sp12_v_b_5')
// (16, 30, 'sp12_v_b_2')
// (16, 31, 'sp12_h_r_1')
// (16, 31, 'sp12_v_b_1')
// (17, 21, 'neigh_op_tnl_1')
// (17, 22, 'neigh_op_lft_1')
// (17, 23, 'neigh_op_bnl_1')
// (17, 31, 'sp12_h_r_2')
// (18, 31, 'sp12_h_r_5')
// (19, 31, 'sp12_h_r_6')
// (20, 31, 'sp12_h_r_9')
// (21, 31, 'sp12_h_r_10')
// (22, 31, 'sp12_h_r_13')
// (23, 31, 'sp12_h_r_14')
// (24, 31, 'sp12_h_r_17')
// (25, 31, 'sp12_h_r_18')
// (26, 31, 'sp12_h_r_21')
// (26, 31, 'sp4_h_r_10')
// (27, 31, 'sp12_h_r_22')
// (27, 31, 'sp4_h_r_23')
// (28, 31, 'sp12_h_l_22')
// (28, 31, 'sp4_h_r_34')
// (29, 31, 'sp4_h_r_47')
// (30, 31, 'sp4_h_l_47')
// (30, 31, 'sp4_h_r_1')
// (31, 31, 'sp4_h_r_12')
// (32, 31, 'sp4_h_r_25')
// (33, 27, 'span4_vert_t_12')
// (33, 28, 'span4_vert_b_12')
// (33, 29, 'span4_vert_b_8')
// (33, 30, 'io_1/D_OUT_0')
// (33, 30, 'io_1/PAD')
// (33, 30, 'local_g1_4')
// (33, 30, 'span4_vert_b_4')
// (33, 31, 'span4_horz_25')
// (33, 31, 'span4_vert_b_0')

reg io_33_31_0 = 0;
// (15, 21, 'neigh_op_tnr_2')
// (15, 22, 'neigh_op_rgt_2')
// (15, 23, 'neigh_op_bnr_2')
// (16, 20, 'sp4_r_v_b_45')
// (16, 21, 'neigh_op_top_2')
// (16, 21, 'sp4_r_v_b_32')
// (16, 22, 'lutff_2/out')
// (16, 22, 'sp4_r_v_b_21')
// (16, 23, 'neigh_op_bot_2')
// (16, 23, 'sp4_r_v_b_8')
// (16, 24, 'sp4_r_v_b_46')
// (16, 25, 'sp4_r_v_b_35')
// (16, 26, 'sp4_r_v_b_22')
// (16, 27, 'sp4_r_v_b_11')
// (16, 28, 'sp4_r_v_b_46')
// (16, 29, 'sp4_r_v_b_35')
// (16, 30, 'sp4_r_v_b_22')
// (16, 31, 'sp4_r_v_b_11')
// (17, 19, 'sp4_v_t_45')
// (17, 20, 'sp4_v_b_45')
// (17, 21, 'neigh_op_tnl_2')
// (17, 21, 'sp4_v_b_32')
// (17, 22, 'neigh_op_lft_2')
// (17, 22, 'sp4_v_b_21')
// (17, 23, 'neigh_op_bnl_2')
// (17, 23, 'sp4_v_b_8')
// (17, 23, 'sp4_v_t_46')
// (17, 24, 'sp4_v_b_46')
// (17, 25, 'sp4_v_b_35')
// (17, 26, 'sp4_v_b_22')
// (17, 27, 'sp4_v_b_11')
// (17, 27, 'sp4_v_t_46')
// (17, 28, 'sp4_v_b_46')
// (17, 29, 'sp4_v_b_35')
// (17, 30, 'sp4_v_b_22')
// (17, 31, 'sp4_h_r_11')
// (17, 31, 'sp4_v_b_11')
// (18, 31, 'sp4_h_r_22')
// (19, 31, 'sp4_h_r_35')
// (20, 31, 'sp4_h_r_46')
// (21, 31, 'sp4_h_l_46')
// (21, 31, 'sp4_h_r_2')
// (22, 31, 'sp4_h_r_15')
// (23, 31, 'sp4_h_r_26')
// (24, 31, 'sp4_h_r_39')
// (25, 31, 'sp4_h_l_39')
// (25, 31, 'sp4_h_r_5')
// (26, 31, 'sp4_h_r_16')
// (27, 31, 'sp4_h_r_29')
// (28, 31, 'sp4_h_r_40')
// (29, 31, 'sp4_h_l_40')
// (29, 31, 'sp4_h_r_1')
// (30, 31, 'sp4_h_r_12')
// (31, 31, 'sp4_h_r_25')
// (32, 31, 'sp4_h_r_36')
// (33, 31, 'io_0/D_OUT_0')
// (33, 31, 'io_0/PAD')
// (33, 31, 'local_g0_4')
// (33, 31, 'span4_horz_36')

wire n1010;
// (15, 21, 'neigh_op_tnr_4')
// (15, 22, 'neigh_op_rgt_4')
// (15, 22, 'sp4_r_v_b_40')
// (15, 22, 'sp4_r_v_b_47')
// (15, 23, 'neigh_op_bnr_4')
// (15, 23, 'sp4_r_v_b_29')
// (15, 23, 'sp4_r_v_b_34')
// (15, 23, 'sp4_r_v_b_39')
// (15, 24, 'sp4_r_v_b_16')
// (15, 24, 'sp4_r_v_b_23')
// (15, 24, 'sp4_r_v_b_26')
// (15, 25, 'sp4_r_v_b_10')
// (15, 25, 'sp4_r_v_b_15')
// (15, 25, 'sp4_r_v_b_5')
// (15, 26, 'sp4_r_v_b_2')
// (16, 21, 'neigh_op_top_4')
// (16, 21, 'sp4_h_r_10')
// (16, 21, 'sp4_v_t_40')
// (16, 21, 'sp4_v_t_47')
// (16, 22, 'lutff_4/out')
// (16, 22, 'sp4_h_r_8')
// (16, 22, 'sp4_v_b_40')
// (16, 22, 'sp4_v_b_47')
// (16, 22, 'sp4_v_t_39')
// (16, 23, 'local_g2_2')
// (16, 23, 'lutff_global/cen')
// (16, 23, 'neigh_op_bot_4')
// (16, 23, 'sp4_v_b_29')
// (16, 23, 'sp4_v_b_34')
// (16, 23, 'sp4_v_b_39')
// (16, 24, 'local_g2_2')
// (16, 24, 'lutff_global/cen')
// (16, 24, 'sp4_v_b_16')
// (16, 24, 'sp4_v_b_23')
// (16, 24, 'sp4_v_b_26')
// (16, 25, 'sp4_v_b_10')
// (16, 25, 'sp4_v_b_15')
// (16, 25, 'sp4_v_b_5')
// (16, 26, 'sp4_v_b_2')
// (17, 21, 'neigh_op_tnl_4')
// (17, 21, 'sp4_h_r_23')
// (17, 22, 'neigh_op_lft_4')
// (17, 22, 'sp4_h_r_21')
// (17, 23, 'neigh_op_bnl_4')
// (18, 21, 'sp4_h_r_34')
// (18, 22, 'sp4_h_r_32')
// (19, 21, 'sp4_h_r_47')
// (19, 22, 'sp4_h_r_45')
// (20, 21, 'sp4_h_l_47')
// (20, 22, 'sp4_h_l_45')
// (20, 22, 'sp4_h_r_11')
// (21, 22, 'sp4_h_r_22')
// (22, 22, 'local_g3_3')
// (22, 22, 'lutff_global/cen')
// (22, 22, 'sp4_h_r_35')
// (23, 22, 'sp4_h_r_46')
// (24, 22, 'sp4_h_l_46')

wire n1011;
// (15, 21, 'sp12_h_r_0')
// (16, 21, 'sp12_h_r_3')
// (17, 21, 'sp12_h_r_4')
// (18, 21, 'sp12_h_r_7')
// (19, 21, 'local_g0_0')
// (19, 21, 'lutff_0/in_0')
// (19, 21, 'sp12_h_r_8')
// (20, 21, 'sp12_h_r_11')
// (21, 21, 'sp12_h_r_12')
// (22, 21, 'sp12_h_r_15')
// (23, 21, 'sp12_h_r_16')
// (24, 21, 'sp12_h_r_19')
// (25, 21, 'sp12_h_r_20')
// (26, 21, 'sp12_h_r_23')
// (26, 32, 'neigh_op_tnr_0')
// (26, 32, 'neigh_op_tnr_4')
// (27, 21, 'sp12_h_l_23')
// (27, 21, 'sp12_v_t_23')
// (27, 22, 'sp12_v_b_23')
// (27, 23, 'sp12_v_b_20')
// (27, 24, 'sp12_v_b_19')
// (27, 25, 'sp12_v_b_16')
// (27, 26, 'sp12_v_b_15')
// (27, 27, 'sp12_v_b_12')
// (27, 28, 'sp12_v_b_11')
// (27, 29, 'sp12_v_b_8')
// (27, 30, 'sp12_v_b_7')
// (27, 31, 'sp12_v_b_4')
// (27, 32, 'neigh_op_top_0')
// (27, 32, 'neigh_op_top_4')
// (27, 32, 'sp12_v_b_3')
// (27, 33, 'io_0/D_IN_0')
// (27, 33, 'span12_vert_0')
// (28, 32, 'neigh_op_tnl_0')
// (28, 32, 'neigh_op_tnl_4')

wire n1012;
// (15, 21, 'sp4_h_r_6')
// (16, 21, 'sp4_h_r_19')
// (17, 21, 'sp4_h_r_30')
// (18, 18, 'sp4_r_v_b_36')
// (18, 19, 'neigh_op_tnr_6')
// (18, 19, 'sp4_r_v_b_25')
// (18, 20, 'neigh_op_rgt_6')
// (18, 20, 'sp4_r_v_b_12')
// (18, 21, 'neigh_op_bnr_6')
// (18, 21, 'sp4_h_r_43')
// (18, 21, 'sp4_r_v_b_1')
// (18, 22, 'sp4_r_v_b_43')
// (18, 23, 'sp4_r_v_b_30')
// (18, 24, 'local_g3_3')
// (18, 24, 'lutff_global/cen')
// (18, 24, 'sp4_r_v_b_19')
// (18, 25, 'sp4_r_v_b_6')
// (19, 14, 'sp12_v_t_23')
// (19, 15, 'sp12_v_b_23')
// (19, 16, 'sp12_v_b_20')
// (19, 17, 'sp12_v_b_19')
// (19, 17, 'sp4_v_t_36')
// (19, 18, 'sp12_v_b_16')
// (19, 18, 'sp4_v_b_36')
// (19, 19, 'neigh_op_top_6')
// (19, 19, 'sp12_v_b_15')
// (19, 19, 'sp4_v_b_25')
// (19, 20, 'lutff_6/out')
// (19, 20, 'sp12_v_b_12')
// (19, 20, 'sp4_v_b_12')
// (19, 21, 'neigh_op_bot_6')
// (19, 21, 'sp12_v_b_11')
// (19, 21, 'sp4_h_l_43')
// (19, 21, 'sp4_h_r_6')
// (19, 21, 'sp4_v_b_1')
// (19, 21, 'sp4_v_t_43')
// (19, 22, 'sp12_v_b_8')
// (19, 22, 'sp4_v_b_43')
// (19, 23, 'sp12_v_b_7')
// (19, 23, 'sp4_v_b_30')
// (19, 24, 'sp12_v_b_4')
// (19, 24, 'sp4_v_b_19')
// (19, 25, 'local_g3_3')
// (19, 25, 'lutff_global/cen')
// (19, 25, 'sp12_v_b_3')
// (19, 25, 'sp4_v_b_6')
// (19, 26, 'sp12_v_b_0')
// (20, 19, 'neigh_op_tnl_6')
// (20, 20, 'neigh_op_lft_6')
// (20, 21, 'local_g1_3')
// (20, 21, 'lutff_global/cen')
// (20, 21, 'neigh_op_bnl_6')
// (20, 21, 'sp4_h_r_19')
// (21, 21, 'sp4_h_r_30')
// (22, 21, 'sp4_h_r_43')
// (23, 21, 'sp4_h_l_43')

wire n1013;
// (15, 22, 'lutff_7/cout')
// (15, 23, 'carry_in')
// (15, 23, 'carry_in_mux')
// (15, 23, 'lutff_0/in_3')

reg n1014 = 0;
// (15, 22, 'neigh_op_tnr_0')
// (15, 23, 'neigh_op_rgt_0')
// (15, 24, 'neigh_op_bnr_0')
// (16, 19, 'sp12_v_t_23')
// (16, 20, 'sp12_v_b_23')
// (16, 21, 'sp12_v_b_20')
// (16, 22, 'neigh_op_top_0')
// (16, 22, 'sp12_v_b_19')
// (16, 23, 'lutff_0/out')
// (16, 23, 'sp12_v_b_16')
// (16, 24, 'neigh_op_bot_0')
// (16, 24, 'sp12_v_b_15')
// (16, 25, 'sp12_v_b_12')
// (16, 26, 'sp12_v_b_11')
// (16, 27, 'sp12_v_b_8')
// (16, 28, 'sp12_v_b_7')
// (16, 29, 'sp12_v_b_4')
// (16, 30, 'sp12_v_b_3')
// (16, 31, 'sp12_h_r_0')
// (16, 31, 'sp12_v_b_0')
// (17, 22, 'neigh_op_tnl_0')
// (17, 23, 'neigh_op_lft_0')
// (17, 24, 'neigh_op_bnl_0')
// (17, 31, 'sp12_h_r_3')
// (18, 31, 'sp12_h_r_4')
// (19, 31, 'sp12_h_r_7')
// (20, 31, 'sp12_h_r_8')
// (21, 31, 'sp12_h_r_11')
// (22, 31, 'sp12_h_r_12')
// (23, 31, 'sp12_h_r_15')
// (23, 31, 'sp4_h_r_9')
// (24, 31, 'sp12_h_r_16')
// (24, 31, 'sp4_h_r_20')
// (25, 31, 'sp12_h_r_19')
// (25, 31, 'sp4_h_r_33')
// (26, 31, 'sp12_h_r_20')
// (26, 31, 'sp4_h_r_44')
// (26, 32, 'sp4_r_v_b_44')
// (27, 31, 'sp12_h_r_23')
// (27, 31, 'sp4_h_l_44')
// (27, 31, 'sp4_v_t_44')
// (27, 32, 'sp4_v_b_44')
// (27, 33, 'io_0/D_OUT_0')
// (27, 33, 'local_g1_1')
// (27, 33, 'span4_vert_33')
// (28, 31, 'sp12_h_l_23')

reg n1015 = 0;
// (15, 22, 'neigh_op_tnr_1')
// (15, 23, 'neigh_op_rgt_1')
// (15, 24, 'neigh_op_bnr_1')
// (16, 20, 'sp12_v_t_22')
// (16, 21, 'sp12_v_b_22')
// (16, 22, 'neigh_op_top_1')
// (16, 22, 'sp12_v_b_21')
// (16, 23, 'lutff_1/out')
// (16, 23, 'sp12_v_b_18')
// (16, 24, 'neigh_op_bot_1')
// (16, 24, 'sp12_v_b_17')
// (16, 25, 'sp12_v_b_14')
// (16, 26, 'sp12_v_b_13')
// (16, 27, 'sp12_v_b_10')
// (16, 28, 'sp12_v_b_9')
// (16, 29, 'sp12_v_b_6')
// (16, 30, 'sp12_v_b_5')
// (16, 31, 'sp12_v_b_2')
// (16, 32, 'sp12_h_r_1')
// (16, 32, 'sp12_v_b_1')
// (17, 22, 'neigh_op_tnl_1')
// (17, 23, 'neigh_op_lft_1')
// (17, 24, 'neigh_op_bnl_1')
// (17, 32, 'sp12_h_r_2')
// (18, 32, 'sp12_h_r_5')
// (19, 32, 'sp12_h_r_6')
// (20, 32, 'sp12_h_r_9')
// (21, 32, 'sp12_h_r_10')
// (22, 32, 'sp12_h_r_13')
// (23, 32, 'sp12_h_r_14')
// (24, 32, 'sp12_h_r_17')
// (25, 32, 'sp12_h_r_18')
// (26, 32, 'sp12_h_r_21')
// (27, 32, 'sp12_h_r_22')
// (28, 32, 'sp12_h_l_22')
// (28, 32, 'sp12_v_t_22')
// (28, 33, 'io_1/D_OUT_0')
// (28, 33, 'local_g1_6')
// (28, 33, 'span12_vert_22')

reg n1016 = 0;
// (15, 22, 'neigh_op_tnr_2')
// (15, 23, 'neigh_op_rgt_2')
// (15, 24, 'neigh_op_bnr_2')
// (16, 9, 'sp12_h_r_0')
// (16, 9, 'sp12_v_t_23')
// (16, 10, 'sp12_v_b_23')
// (16, 11, 'sp12_v_b_20')
// (16, 12, 'sp12_v_b_19')
// (16, 13, 'sp12_v_b_16')
// (16, 14, 'sp12_v_b_15')
// (16, 15, 'sp12_v_b_12')
// (16, 16, 'sp12_v_b_11')
// (16, 17, 'sp12_v_b_8')
// (16, 18, 'sp12_v_b_7')
// (16, 19, 'sp12_v_b_4')
// (16, 20, 'sp12_v_b_3')
// (16, 21, 'sp12_v_b_0')
// (16, 21, 'sp12_v_t_23')
// (16, 22, 'neigh_op_top_2')
// (16, 22, 'sp12_v_b_23')
// (16, 23, 'lutff_2/out')
// (16, 23, 'sp12_v_b_20')
// (16, 24, 'neigh_op_bot_2')
// (16, 24, 'sp12_v_b_19')
// (16, 25, 'sp12_v_b_16')
// (16, 26, 'sp12_v_b_15')
// (16, 27, 'sp12_v_b_12')
// (16, 28, 'sp12_v_b_11')
// (16, 29, 'sp12_v_b_8')
// (16, 30, 'sp12_v_b_7')
// (16, 31, 'sp12_v_b_4')
// (16, 32, 'sp12_v_b_3')
// (16, 33, 'span12_vert_0')
// (17, 9, 'sp12_h_r_3')
// (17, 22, 'neigh_op_tnl_2')
// (17, 23, 'neigh_op_lft_2')
// (17, 24, 'neigh_op_bnl_2')
// (18, 9, 'sp12_h_r_4')
// (19, 9, 'sp12_h_r_7')
// (20, 9, 'sp12_h_r_8')
// (21, 9, 'sp12_h_r_11')
// (21, 9, 'sp4_h_r_7')
// (22, 9, 'sp12_h_r_12')
// (22, 9, 'sp4_h_r_18')
// (23, 9, 'sp12_h_r_15')
// (23, 9, 'sp4_h_r_31')
// (24, 9, 'sp12_h_r_16')
// (24, 9, 'sp4_h_r_42')
// (25, 9, 'sp12_h_r_19')
// (25, 9, 'sp4_h_l_42')
// (25, 9, 'sp4_h_r_7')
// (26, 9, 'sp12_h_r_20')
// (26, 9, 'sp4_h_r_18')
// (27, 9, 'sp12_h_r_23')
// (27, 9, 'sp4_h_r_31')
// (28, 6, 'sp4_r_v_b_42')
// (28, 7, 'sp4_r_v_b_31')
// (28, 8, 'sp4_r_v_b_18')
// (28, 9, 'sp12_h_l_23')
// (28, 9, 'sp4_h_r_42')
// (28, 9, 'sp4_r_v_b_7')
// (29, 5, 'sp4_h_r_0')
// (29, 5, 'sp4_v_t_42')
// (29, 6, 'sp4_v_b_42')
// (29, 7, 'sp4_v_b_31')
// (29, 8, 'sp4_v_b_18')
// (29, 9, 'sp4_h_l_42')
// (29, 9, 'sp4_v_b_7')
// (30, 5, 'sp4_h_r_13')
// (31, 5, 'sp4_h_r_24')
// (32, 5, 'sp4_h_r_37')
// (33, 1, 'span4_vert_t_14')
// (33, 2, 'io_1/D_OUT_0')
// (33, 2, 'local_g1_6')
// (33, 2, 'span4_vert_b_14')
// (33, 3, 'span4_vert_b_10')
// (33, 4, 'span4_vert_b_6')
// (33, 5, 'span4_horz_37')
// (33, 5, 'span4_vert_b_2')

reg n1017 = 0;
// (15, 22, 'neigh_op_tnr_3')
// (15, 23, 'neigh_op_rgt_3')
// (15, 24, 'neigh_op_bnr_3')
// (16, 22, 'neigh_op_top_3')
// (16, 22, 'sp12_h_r_1')
// (16, 22, 'sp12_v_t_22')
// (16, 23, 'lutff_3/out')
// (16, 23, 'sp12_v_b_22')
// (16, 24, 'neigh_op_bot_3')
// (16, 24, 'sp12_v_b_21')
// (16, 25, 'sp12_v_b_18')
// (16, 26, 'sp12_v_b_17')
// (16, 27, 'sp12_v_b_14')
// (16, 28, 'sp12_v_b_13')
// (16, 29, 'sp12_v_b_10')
// (16, 30, 'sp12_v_b_9')
// (16, 31, 'sp12_v_b_6')
// (16, 32, 'sp12_v_b_5')
// (16, 33, 'span12_vert_2')
// (17, 22, 'neigh_op_tnl_3')
// (17, 22, 'sp12_h_r_2')
// (17, 23, 'neigh_op_lft_3')
// (17, 24, 'neigh_op_bnl_3')
// (18, 22, 'sp12_h_r_5')
// (19, 22, 'sp12_h_r_6')
// (20, 22, 'sp12_h_r_9')
// (21, 22, 'sp12_h_r_10')
// (22, 22, 'sp12_h_r_13')
// (23, 22, 'sp12_h_r_14')
// (24, 22, 'sp12_h_r_17')
// (25, 22, 'sp12_h_r_18')
// (26, 22, 'sp12_h_r_21')
// (26, 22, 'sp4_h_r_10')
// (27, 22, 'sp12_h_r_22')
// (27, 22, 'sp4_h_r_23')
// (28, 22, 'sp12_h_l_22')
// (28, 22, 'sp4_h_r_34')
// (29, 15, 'sp4_r_v_b_41')
// (29, 16, 'sp4_r_v_b_28')
// (29, 17, 'sp4_r_v_b_17')
// (29, 18, 'sp4_r_v_b_4')
// (29, 19, 'sp4_r_v_b_41')
// (29, 20, 'sp4_r_v_b_28')
// (29, 21, 'sp4_r_v_b_17')
// (29, 22, 'sp4_h_r_47')
// (29, 22, 'sp4_r_v_b_4')
// (30, 14, 'sp4_h_r_4')
// (30, 14, 'sp4_v_t_41')
// (30, 15, 'sp4_v_b_41')
// (30, 16, 'sp4_v_b_28')
// (30, 17, 'sp4_v_b_17')
// (30, 18, 'sp4_v_b_4')
// (30, 18, 'sp4_v_t_41')
// (30, 19, 'sp4_v_b_41')
// (30, 20, 'sp4_v_b_28')
// (30, 21, 'sp4_v_b_17')
// (30, 22, 'sp4_h_l_47')
// (30, 22, 'sp4_v_b_4')
// (31, 14, 'sp4_h_r_17')
// (32, 14, 'sp4_h_r_28')
// (33, 14, 'io_1/D_OUT_0')
// (33, 14, 'local_g1_4')
// (33, 14, 'span4_horz_28')

reg n1018 = 0;
// (15, 22, 'neigh_op_tnr_4')
// (15, 23, 'neigh_op_rgt_4')
// (15, 24, 'neigh_op_bnr_4')
// (16, 15, 'sp12_v_t_23')
// (16, 16, 'sp12_v_b_23')
// (16, 17, 'sp12_v_b_20')
// (16, 18, 'sp12_v_b_19')
// (16, 19, 'sp12_v_b_16')
// (16, 20, 'sp12_v_b_15')
// (16, 21, 'sp12_v_b_12')
// (16, 22, 'neigh_op_top_4')
// (16, 22, 'sp12_v_b_11')
// (16, 23, 'lutff_4/out')
// (16, 23, 'sp12_v_b_8')
// (16, 24, 'neigh_op_bot_4')
// (16, 24, 'sp12_v_b_7')
// (16, 25, 'sp12_v_b_4')
// (16, 26, 'sp12_v_b_3')
// (16, 27, 'sp12_h_r_0')
// (16, 27, 'sp12_v_b_0')
// (17, 22, 'neigh_op_tnl_4')
// (17, 23, 'neigh_op_lft_4')
// (17, 24, 'neigh_op_bnl_4')
// (17, 27, 'sp12_h_r_3')
// (18, 27, 'sp12_h_r_4')
// (19, 27, 'sp12_h_r_7')
// (20, 27, 'sp12_h_r_8')
// (21, 27, 'sp12_h_r_11')
// (22, 27, 'sp12_h_r_12')
// (23, 27, 'sp12_h_r_15')
// (24, 27, 'sp12_h_r_16')
// (25, 27, 'sp12_h_r_19')
// (26, 27, 'sp12_h_r_20')
// (27, 27, 'sp12_h_r_23')
// (28, 15, 'sp12_h_r_0')
// (28, 15, 'sp12_v_t_23')
// (28, 16, 'sp12_v_b_23')
// (28, 17, 'sp12_v_b_20')
// (28, 18, 'sp12_v_b_19')
// (28, 19, 'sp12_v_b_16')
// (28, 20, 'sp12_v_b_15')
// (28, 21, 'sp12_v_b_12')
// (28, 22, 'sp12_v_b_11')
// (28, 23, 'sp12_v_b_8')
// (28, 24, 'sp12_v_b_7')
// (28, 25, 'sp12_v_b_4')
// (28, 26, 'sp12_v_b_3')
// (28, 27, 'sp12_h_l_23')
// (28, 27, 'sp12_v_b_0')
// (29, 15, 'sp12_h_r_3')
// (30, 15, 'sp12_h_r_4')
// (31, 15, 'sp12_h_r_7')
// (32, 15, 'sp12_h_r_8')
// (33, 15, 'io_0/D_OUT_0')
// (33, 15, 'local_g0_0')
// (33, 15, 'span12_horz_8')

reg n1019 = 0;
// (15, 22, 'neigh_op_tnr_5')
// (15, 23, 'neigh_op_rgt_5')
// (15, 23, 'sp12_h_r_1')
// (15, 24, 'neigh_op_bnr_5')
// (16, 22, 'neigh_op_top_5')
// (16, 23, 'lutff_5/out')
// (16, 23, 'sp12_h_r_2')
// (16, 24, 'neigh_op_bot_5')
// (17, 22, 'neigh_op_tnl_5')
// (17, 23, 'neigh_op_lft_5')
// (17, 23, 'sp12_h_r_5')
// (17, 24, 'neigh_op_bnl_5')
// (18, 23, 'sp12_h_r_6')
// (19, 23, 'sp12_h_r_9')
// (20, 23, 'sp12_h_r_10')
// (21, 23, 'sp12_h_r_13')
// (22, 23, 'sp12_h_r_14')
// (23, 23, 'sp12_h_r_17')
// (24, 23, 'sp12_h_r_18')
// (25, 23, 'sp12_h_r_21')
// (25, 23, 'sp4_h_r_10')
// (26, 23, 'sp12_h_r_22')
// (26, 23, 'sp4_h_r_23')
// (27, 23, 'sp12_h_l_22')
// (27, 23, 'sp4_h_r_34')
// (28, 16, 'sp4_r_v_b_42')
// (28, 17, 'sp4_r_v_b_31')
// (28, 18, 'sp4_r_v_b_18')
// (28, 19, 'sp4_r_v_b_7')
// (28, 20, 'sp4_r_v_b_41')
// (28, 21, 'sp4_r_v_b_28')
// (28, 22, 'sp4_r_v_b_17')
// (28, 23, 'sp4_h_r_47')
// (28, 23, 'sp4_r_v_b_4')
// (29, 15, 'sp4_h_r_7')
// (29, 15, 'sp4_v_t_42')
// (29, 16, 'sp4_v_b_42')
// (29, 17, 'sp4_v_b_31')
// (29, 18, 'sp4_v_b_18')
// (29, 19, 'sp4_v_b_7')
// (29, 19, 'sp4_v_t_41')
// (29, 20, 'sp4_v_b_41')
// (29, 21, 'sp4_v_b_28')
// (29, 22, 'sp4_v_b_17')
// (29, 23, 'sp4_h_l_47')
// (29, 23, 'sp4_v_b_4')
// (30, 15, 'sp4_h_r_18')
// (31, 15, 'sp4_h_r_31')
// (32, 15, 'sp4_h_r_42')
// (33, 15, 'io_1/D_OUT_0')
// (33, 15, 'local_g1_2')
// (33, 15, 'span4_horz_42')

reg n1020 = 0;
// (15, 22, 'neigh_op_tnr_6')
// (15, 23, 'neigh_op_rgt_6')
// (15, 24, 'neigh_op_bnr_6')
// (16, 21, 'sp4_r_v_b_37')
// (16, 22, 'neigh_op_top_6')
// (16, 22, 'sp4_r_v_b_24')
// (16, 23, 'lutff_6/out')
// (16, 23, 'sp4_r_v_b_13')
// (16, 24, 'neigh_op_bot_6')
// (16, 24, 'sp4_r_v_b_0')
// (17, 20, 'sp4_h_r_5')
// (17, 20, 'sp4_v_t_37')
// (17, 21, 'sp4_v_b_37')
// (17, 22, 'neigh_op_tnl_6')
// (17, 22, 'sp4_v_b_24')
// (17, 23, 'neigh_op_lft_6')
// (17, 23, 'sp4_v_b_13')
// (17, 24, 'neigh_op_bnl_6')
// (17, 24, 'sp4_v_b_0')
// (18, 20, 'sp4_h_r_16')
// (19, 20, 'sp4_h_r_29')
// (20, 20, 'sp4_h_r_40')
// (21, 20, 'sp4_h_l_40')
// (21, 20, 'sp4_h_r_5')
// (22, 20, 'sp4_h_r_16')
// (23, 20, 'sp4_h_r_29')
// (24, 20, 'sp4_h_r_40')
// (25, 20, 'sp4_h_l_40')
// (25, 20, 'sp4_h_r_5')
// (26, 20, 'sp4_h_r_16')
// (27, 20, 'sp4_h_r_29')
// (28, 17, 'sp4_r_v_b_46')
// (28, 18, 'sp4_r_v_b_35')
// (28, 19, 'sp4_r_v_b_22')
// (28, 20, 'sp4_h_r_40')
// (28, 20, 'sp4_r_v_b_11')
// (29, 16, 'sp4_h_r_4')
// (29, 16, 'sp4_v_t_46')
// (29, 17, 'sp4_v_b_46')
// (29, 18, 'sp4_v_b_35')
// (29, 19, 'sp4_v_b_22')
// (29, 20, 'sp4_h_l_40')
// (29, 20, 'sp4_v_b_11')
// (30, 16, 'sp4_h_r_17')
// (31, 16, 'sp4_h_r_28')
// (32, 16, 'sp4_h_r_41')
// (33, 16, 'io_0/D_OUT_0')
// (33, 16, 'local_g1_1')
// (33, 16, 'span4_horz_41')

reg n1021 = 0;
// (15, 22, 'sp12_h_r_1')
// (16, 22, 'sp12_h_r_2')
// (17, 21, 'neigh_op_tnr_7')
// (17, 22, 'neigh_op_rgt_7')
// (17, 22, 'sp12_h_r_5')
// (17, 23, 'neigh_op_bnr_7')
// (18, 21, 'neigh_op_top_7')
// (18, 22, 'local_g1_7')
// (18, 22, 'lutff_7/in_1')
// (18, 22, 'lutff_7/out')
// (18, 22, 'sp12_h_r_6')
// (18, 23, 'neigh_op_bot_7')
// (19, 21, 'neigh_op_tnl_7')
// (19, 22, 'neigh_op_lft_7')
// (19, 22, 'sp12_h_r_9')
// (19, 23, 'neigh_op_bnl_7')
// (20, 22, 'sp12_h_r_10')
// (21, 22, 'sp12_h_r_13')
// (22, 22, 'sp12_h_r_14')
// (23, 22, 'sp12_h_r_17')
// (24, 22, 'sp12_h_r_18')
// (25, 22, 'sp12_h_r_21')
// (26, 22, 'sp12_h_r_22')
// (27, 22, 'sp12_h_l_22')
// (27, 22, 'sp12_v_t_22')
// (27, 23, 'sp12_v_b_22')
// (27, 24, 'sp12_v_b_21')
// (27, 25, 'sp12_v_b_18')
// (27, 26, 'sp12_v_b_17')
// (27, 27, 'sp12_v_b_14')
// (27, 28, 'sp12_v_b_13')
// (27, 29, 'sp12_v_b_10')
// (27, 30, 'sp12_v_b_9')
// (27, 31, 'sp12_v_b_6')
// (27, 32, 'sp12_v_b_5')
// (27, 33, 'io_0/OUT_ENB')
// (27, 33, 'local_g1_2')
// (27, 33, 'span12_vert_2')

reg n1022 = 0;
// (15, 23, 'neigh_op_tnr_0')
// (15, 24, 'neigh_op_rgt_0')
// (15, 25, 'neigh_op_bnr_0')
// (16, 20, 'sp12_v_t_23')
// (16, 21, 'sp12_v_b_23')
// (16, 22, 'sp12_v_b_20')
// (16, 23, 'neigh_op_top_0')
// (16, 23, 'sp12_v_b_19')
// (16, 24, 'lutff_0/out')
// (16, 24, 'sp12_v_b_16')
// (16, 25, 'neigh_op_bot_0')
// (16, 25, 'sp12_v_b_15')
// (16, 26, 'sp12_v_b_12')
// (16, 27, 'sp12_v_b_11')
// (16, 28, 'sp12_v_b_8')
// (16, 29, 'sp12_v_b_7')
// (16, 30, 'sp12_v_b_4')
// (16, 31, 'sp12_v_b_3')
// (16, 32, 'sp12_h_r_0')
// (16, 32, 'sp12_v_b_0')
// (17, 23, 'neigh_op_tnl_0')
// (17, 24, 'neigh_op_lft_0')
// (17, 25, 'neigh_op_bnl_0')
// (17, 32, 'sp12_h_r_3')
// (18, 32, 'sp12_h_r_4')
// (19, 32, 'sp12_h_r_7')
// (20, 32, 'sp12_h_r_8')
// (21, 32, 'sp12_h_r_11')
// (22, 32, 'sp12_h_r_12')
// (23, 32, 'sp12_h_r_15')
// (24, 32, 'sp12_h_r_16')
// (25, 32, 'sp12_h_r_19')
// (25, 32, 'sp4_h_r_11')
// (26, 32, 'sp12_h_r_20')
// (26, 32, 'sp4_h_r_22')
// (27, 32, 'sp12_h_r_23')
// (27, 32, 'sp4_h_r_35')
// (28, 32, 'sp12_h_l_23')
// (28, 32, 'sp4_h_r_46')
// (29, 32, 'sp4_h_l_46')
// (29, 32, 'sp4_v_t_41')
// (29, 33, 'io_1/D_OUT_0')
// (29, 33, 'local_g0_1')
// (29, 33, 'span4_vert_41')

reg n1023 = 0;
// (15, 23, 'neigh_op_tnr_2')
// (15, 24, 'neigh_op_rgt_2')
// (15, 25, 'neigh_op_bnr_2')
// (16, 22, 'sp12_h_r_0')
// (16, 22, 'sp12_v_t_23')
// (16, 23, 'neigh_op_top_2')
// (16, 23, 'sp12_v_b_23')
// (16, 24, 'lutff_2/out')
// (16, 24, 'sp12_v_b_20')
// (16, 25, 'neigh_op_bot_2')
// (16, 25, 'sp12_v_b_19')
// (16, 26, 'sp12_v_b_16')
// (16, 27, 'sp12_v_b_15')
// (16, 28, 'sp12_v_b_12')
// (16, 29, 'sp12_v_b_11')
// (16, 30, 'sp12_v_b_8')
// (16, 31, 'sp12_v_b_7')
// (16, 32, 'sp12_v_b_4')
// (16, 33, 'span12_vert_3')
// (17, 22, 'sp12_h_r_3')
// (17, 23, 'neigh_op_tnl_2')
// (17, 24, 'neigh_op_lft_2')
// (17, 25, 'neigh_op_bnl_2')
// (18, 22, 'sp12_h_r_4')
// (19, 22, 'sp12_h_r_7')
// (20, 22, 'sp12_h_r_8')
// (21, 22, 'sp12_h_r_11')
// (22, 22, 'sp12_h_r_12')
// (23, 22, 'sp12_h_r_15')
// (24, 22, 'sp12_h_r_16')
// (25, 22, 'sp12_h_r_19')
// (26, 22, 'sp12_h_r_20')
// (27, 22, 'sp12_h_r_23')
// (27, 27, 'sp4_r_v_b_41')
// (27, 28, 'sp4_r_v_b_28')
// (27, 29, 'sp4_r_v_b_17')
// (27, 30, 'sp4_r_v_b_4')
// (27, 31, 'sp4_r_v_b_37')
// (27, 32, 'sp4_r_v_b_24')
// (28, 22, 'sp12_h_l_23')
// (28, 22, 'sp12_v_t_23')
// (28, 23, 'sp12_v_b_23')
// (28, 24, 'sp12_v_b_20')
// (28, 25, 'sp12_v_b_19')
// (28, 26, 'sp12_v_b_16')
// (28, 26, 'sp4_v_t_41')
// (28, 27, 'sp12_v_b_15')
// (28, 27, 'sp4_v_b_41')
// (28, 28, 'sp12_v_b_12')
// (28, 28, 'sp4_v_b_28')
// (28, 29, 'sp12_v_b_11')
// (28, 29, 'sp4_v_b_17')
// (28, 30, 'sp12_v_b_8')
// (28, 30, 'sp4_v_b_4')
// (28, 30, 'sp4_v_t_37')
// (28, 31, 'sp12_v_b_7')
// (28, 31, 'sp4_v_b_37')
// (28, 32, 'sp12_v_b_4')
// (28, 32, 'sp4_v_b_24')
// (28, 33, 'span12_vert_3')
// (28, 33, 'span4_horz_r_2')
// (28, 33, 'span4_vert_13')
// (29, 33, 'span4_horz_r_6')
// (30, 33, 'io_1/D_OUT_0')
// (30, 33, 'local_g1_2')
// (30, 33, 'span4_horz_r_10')
// (31, 33, 'span4_horz_r_14')
// (32, 33, 'span4_horz_l_14')

reg n1024 = 0;
// (15, 23, 'sp12_h_r_0')
// (16, 23, 'sp12_h_r_3')
// (17, 23, 'sp12_h_r_4')
// (18, 22, 'neigh_op_tnr_0')
// (18, 23, 'neigh_op_rgt_0')
// (18, 23, 'sp12_h_r_7')
// (18, 24, 'neigh_op_bnr_0')
// (19, 22, 'neigh_op_top_0')
// (19, 23, 'local_g0_0')
// (19, 23, 'lutff_0/in_0')
// (19, 23, 'lutff_0/out')
// (19, 23, 'sp12_h_r_8')
// (19, 24, 'neigh_op_bot_0')
// (20, 22, 'neigh_op_tnl_0')
// (20, 23, 'neigh_op_lft_0')
// (20, 23, 'sp12_h_r_11')
// (20, 24, 'neigh_op_bnl_0')
// (21, 23, 'sp12_h_r_12')
// (22, 23, 'sp12_h_r_15')
// (23, 23, 'sp12_h_r_16')
// (24, 23, 'sp12_h_r_19')
// (25, 23, 'sp12_h_r_20')
// (26, 23, 'sp12_h_r_23')
// (26, 28, 'sp4_r_v_b_41')
// (26, 29, 'sp4_r_v_b_28')
// (26, 30, 'sp4_r_v_b_17')
// (26, 31, 'sp4_r_v_b_4')
// (26, 32, 'sp4_r_v_b_42')
// (27, 23, 'sp12_h_l_23')
// (27, 23, 'sp12_v_t_23')
// (27, 24, 'sp12_v_b_23')
// (27, 25, 'sp12_v_b_20')
// (27, 26, 'sp12_v_b_19')
// (27, 27, 'sp12_v_b_16')
// (27, 27, 'sp4_v_t_41')
// (27, 28, 'sp12_v_b_15')
// (27, 28, 'sp4_v_b_41')
// (27, 29, 'sp12_v_b_12')
// (27, 29, 'sp4_v_b_28')
// (27, 30, 'sp12_v_b_11')
// (27, 30, 'sp4_v_b_17')
// (27, 31, 'sp12_v_b_8')
// (27, 31, 'sp4_v_b_4')
// (27, 31, 'sp4_v_t_42')
// (27, 32, 'sp12_v_b_7')
// (27, 32, 'sp4_v_b_42')
// (27, 33, 'span12_vert_4')
// (27, 33, 'span4_horz_r_1')
// (27, 33, 'span4_vert_31')
// (28, 33, 'span4_horz_r_5')
// (29, 33, 'span4_horz_r_9')
// (30, 33, 'io_1/OUT_ENB')
// (30, 33, 'local_g1_5')
// (30, 33, 'span4_horz_r_13')
// (31, 33, 'span4_horz_l_13')

wire n1025;
// (15, 23, 'sp4_h_r_1')
// (16, 19, 'sp4_r_v_b_44')
// (16, 20, 'local_g2_1')
// (16, 20, 'lutff_0/in_3')
// (16, 20, 'sp4_r_v_b_33')
// (16, 21, 'sp4_r_v_b_20')
// (16, 22, 'sp4_r_v_b_9')
// (16, 23, 'sp4_h_r_12')
// (17, 18, 'sp4_v_t_44')
// (17, 19, 'sp4_v_b_44')
// (17, 20, 'sp4_v_b_33')
// (17, 21, 'neigh_op_tnr_2')
// (17, 21, 'sp4_v_b_20')
// (17, 22, 'neigh_op_rgt_2')
// (17, 22, 'sp4_h_r_9')
// (17, 22, 'sp4_v_b_9')
// (17, 23, 'neigh_op_bnr_2')
// (17, 23, 'sp4_h_r_25')
// (18, 20, 'sp12_v_t_23')
// (18, 20, 'sp4_r_v_b_45')
// (18, 21, 'neigh_op_top_2')
// (18, 21, 'sp12_v_b_23')
// (18, 21, 'sp4_r_v_b_32')
// (18, 22, 'local_g3_2')
// (18, 22, 'lutff_0/in_3')
// (18, 22, 'lutff_2/out')
// (18, 22, 'lutff_4/in_3')
// (18, 22, 'lutff_5/in_0')
// (18, 22, 'lutff_6/in_3')
// (18, 22, 'lutff_7/in_0')
// (18, 22, 'sp12_v_b_20')
// (18, 22, 'sp4_h_r_20')
// (18, 22, 'sp4_r_v_b_21')
// (18, 23, 'neigh_op_bot_2')
// (18, 23, 'sp12_v_b_19')
// (18, 23, 'sp4_h_r_36')
// (18, 23, 'sp4_r_v_b_8')
// (18, 24, 'sp12_v_b_16')
// (18, 24, 'sp4_r_v_b_43')
// (18, 25, 'sp12_v_b_15')
// (18, 25, 'sp4_r_v_b_30')
// (18, 26, 'local_g3_4')
// (18, 26, 'lutff_0/in_3')
// (18, 26, 'sp12_v_b_12')
// (18, 26, 'sp4_r_v_b_19')
// (18, 27, 'sp12_v_b_11')
// (18, 27, 'sp4_r_v_b_6')
// (18, 28, 'sp12_v_b_8')
// (18, 29, 'sp12_v_b_7')
// (18, 30, 'sp12_v_b_4')
// (18, 31, 'sp12_v_b_3')
// (18, 32, 'sp12_v_b_0')
// (19, 19, 'sp4_v_t_45')
// (19, 20, 'local_g2_5')
// (19, 20, 'lutff_0/in_3')
// (19, 20, 'lutff_1/in_0')
// (19, 20, 'lutff_2/in_3')
// (19, 20, 'lutff_3/in_0')
// (19, 20, 'lutff_4/in_3')
// (19, 20, 'sp4_v_b_45')
// (19, 21, 'local_g3_2')
// (19, 21, 'lutff_0/in_3')
// (19, 21, 'lutff_1/in_0')
// (19, 21, 'lutff_2/in_3')
// (19, 21, 'lutff_3/in_0')
// (19, 21, 'lutff_4/in_3')
// (19, 21, 'lutff_5/in_0')
// (19, 21, 'lutff_6/in_3')
// (19, 21, 'lutff_7/in_0')
// (19, 21, 'neigh_op_tnl_2')
// (19, 21, 'sp4_v_b_32')
// (19, 22, 'neigh_op_lft_2')
// (19, 22, 'sp4_h_r_33')
// (19, 22, 'sp4_v_b_21')
// (19, 23, 'local_g3_2')
// (19, 23, 'lutff_0/in_3')
// (19, 23, 'lutff_1/in_0')
// (19, 23, 'lutff_2/in_3')
// (19, 23, 'lutff_3/in_0')
// (19, 23, 'lutff_4/in_3')
// (19, 23, 'lutff_5/in_0')
// (19, 23, 'lutff_6/in_3')
// (19, 23, 'lutff_7/in_0')
// (19, 23, 'neigh_op_bnl_2')
// (19, 23, 'sp4_h_l_36')
// (19, 23, 'sp4_v_b_8')
// (19, 23, 'sp4_v_t_43')
// (19, 24, 'local_g3_3')
// (19, 24, 'lutff_global/cen')
// (19, 24, 'sp4_v_b_43')
// (19, 25, 'sp4_v_b_30')
// (19, 26, 'sp4_v_b_19')
// (19, 27, 'sp4_v_b_6')
// (20, 22, 'local_g3_4')
// (20, 22, 'lutff_2/in_3')
// (20, 22, 'sp4_h_r_44')
// (21, 22, 'sp4_h_l_44')
// (21, 22, 'sp4_h_r_5')
// (22, 22, 'sp4_h_r_16')
// (23, 22, 'sp4_h_r_29')
// (24, 22, 'local_g3_0')
// (24, 22, 'lutff_4/in_3')
// (24, 22, 'sp4_h_r_40')
// (25, 22, 'sp4_h_l_40')

wire n1026;
// (15, 24, 'carry_in_mux')
// (15, 24, 'lutff_0/in_3')

wire n1027;
// (15, 24, 'lutff_0/cout')
// (15, 24, 'lutff_1/in_3')

wire n1028;
// (15, 24, 'lutff_1/cout')
// (15, 24, 'lutff_2/in_3')

wire n1029;
// (15, 24, 'lutff_2/cout')
// (15, 24, 'lutff_3/in_3')

wire n1030;
// (15, 24, 'lutff_3/cout')
// (15, 24, 'lutff_4/in_3')

wire n1031;
// (15, 24, 'lutff_4/cout')
// (15, 24, 'lutff_5/in_3')

wire n1032;
// (15, 24, 'lutff_5/cout')
// (15, 24, 'lutff_6/in_3')

wire n1033;
// (15, 24, 'lutff_6/cout')
// (15, 24, 'lutff_7/in_3')

wire n1034;
// (15, 24, 'lutff_7/cout')
// (15, 25, 'carry_in')
// (15, 25, 'carry_in_mux')
// (15, 25, 'lutff_0/in_3')

reg n1035 = 0;
// (15, 24, 'sp4_h_r_3')
// (16, 24, 'sp4_h_r_14')
// (17, 24, 'sp4_h_r_27')
// (18, 24, 'local_g2_6')
// (18, 24, 'lutff_1/in_3')
// (18, 24, 'sp4_h_r_38')
// (19, 24, 'sp4_h_l_38')
// (19, 24, 'sp4_h_r_7')
// (20, 24, 'sp4_h_r_18')
// (21, 24, 'sp4_h_r_31')
// (22, 21, 'neigh_op_tnr_5')
// (22, 21, 'sp4_r_v_b_39')
// (22, 22, 'neigh_op_rgt_5')
// (22, 22, 'sp4_r_v_b_26')
// (22, 23, 'neigh_op_bnr_5')
// (22, 23, 'sp4_r_v_b_15')
// (22, 24, 'sp4_h_r_42')
// (22, 24, 'sp4_r_v_b_2')
// (23, 20, 'sp4_v_t_39')
// (23, 21, 'neigh_op_top_5')
// (23, 21, 'sp4_v_b_39')
// (23, 22, 'lutff_5/out')
// (23, 22, 'sp4_v_b_26')
// (23, 23, 'neigh_op_bot_5')
// (23, 23, 'sp4_v_b_15')
// (23, 24, 'sp4_h_l_42')
// (23, 24, 'sp4_v_b_2')
// (24, 21, 'neigh_op_tnl_5')
// (24, 22, 'neigh_op_lft_5')
// (24, 23, 'neigh_op_bnl_5')

wire n1036;
// (15, 25, 'lutff_0/cout')
// (15, 25, 'lutff_1/in_3')

wire n1037;
// (15, 25, 'lutff_1/cout')
// (15, 25, 'lutff_2/in_3')

wire n1038;
// (15, 25, 'lutff_2/cout')
// (15, 25, 'lutff_3/in_3')

wire n1039;
// (15, 25, 'lutff_3/cout')
// (15, 25, 'lutff_4/in_3')

wire n1040;
// (15, 25, 'lutff_4/cout')
// (15, 25, 'lutff_5/in_3')

wire n1041;
// (15, 25, 'lutff_5/cout')
// (15, 25, 'lutff_6/in_3')

wire n1042;
// (15, 25, 'lutff_6/cout')
// (15, 25, 'lutff_7/in_3')

wire n1043;
// (15, 25, 'lutff_7/cout')
// (15, 26, 'carry_in')
// (15, 26, 'carry_in_mux')
// (15, 26, 'lutff_0/in_3')

reg n1044 = 0;
// (15, 25, 'neigh_op_tnr_5')
// (15, 26, 'neigh_op_rgt_5')
// (15, 27, 'neigh_op_bnr_5')
// (16, 25, 'neigh_op_top_5')
// (16, 26, 'lutff_5/out')
// (16, 27, 'neigh_op_bot_5')
// (17, 25, 'local_g3_5')
// (17, 25, 'lutff_3/in_3')
// (17, 25, 'neigh_op_tnl_5')
// (17, 26, 'neigh_op_lft_5')
// (17, 27, 'neigh_op_bnl_5')

wire n1045;
// (15, 26, 'lutff_0/cout')
// (15, 26, 'lutff_1/in_3')

wire n1046;
// (15, 26, 'lutff_1/cout')
// (15, 26, 'lutff_2/in_3')

reg n1047 = 0;
// (16, 6, 'sp12_v_t_23')
// (16, 7, 'sp12_v_b_23')
// (16, 8, 'sp12_v_b_20')
// (16, 9, 'sp12_v_b_19')
// (16, 10, 'local_g2_0')
// (16, 10, 'lutff_5/in_3')
// (16, 10, 'sp12_v_b_16')
// (16, 11, 'sp12_v_b_15')
// (16, 12, 'sp12_v_b_12')
// (16, 13, 'sp12_v_b_11')
// (16, 14, 'sp12_v_b_8')
// (16, 15, 'sp12_v_b_7')
// (16, 16, 'sp12_v_b_4')
// (16, 17, 'sp12_v_b_3')
// (16, 18, 'sp12_h_r_0')
// (16, 18, 'sp12_v_b_0')
// (17, 18, 'sp12_h_r_3')
// (18, 18, 'sp12_h_r_4')
// (19, 18, 'sp12_h_r_7')
// (20, 18, 'sp12_h_r_8')
// (21, 17, 'neigh_op_tnr_2')
// (21, 18, 'neigh_op_rgt_2')
// (21, 18, 'sp12_h_r_11')
// (21, 19, 'neigh_op_bnr_2')
// (22, 17, 'neigh_op_top_2')
// (22, 18, 'lutff_2/out')
// (22, 18, 'sp12_h_r_12')
// (22, 19, 'neigh_op_bot_2')
// (23, 17, 'neigh_op_tnl_2')
// (23, 18, 'neigh_op_lft_2')
// (23, 18, 'sp12_h_r_15')
// (23, 19, 'neigh_op_bnl_2')
// (24, 18, 'sp12_h_r_16')
// (25, 18, 'sp12_h_r_19')
// (26, 18, 'sp12_h_r_20')
// (27, 18, 'sp12_h_r_23')
// (28, 18, 'sp12_h_l_23')

wire n1048;
// (16, 7, 'lutff_0/cout')
// (16, 7, 'lutff_1/in_3')

wire n1049;
// (16, 7, 'lutff_1/cout')
// (16, 7, 'lutff_2/in_3')

wire n1050;
// (16, 7, 'lutff_2/cout')
// (16, 7, 'lutff_3/in_3')

wire n1051;
// (16, 7, 'lutff_3/cout')
// (16, 7, 'lutff_4/in_3')

wire n1052;
// (16, 7, 'lutff_4/cout')
// (16, 7, 'lutff_5/in_3')

reg n1053 = 0;
// (16, 7, 'sp4_r_v_b_44')
// (16, 8, 'sp4_r_v_b_33')
// (16, 9, 'sp4_r_v_b_20')
// (16, 10, 'sp4_r_v_b_9')
// (16, 11, 'sp4_r_v_b_43')
// (16, 12, 'sp4_r_v_b_30')
// (16, 13, 'sp4_r_v_b_19')
// (16, 14, 'sp4_r_v_b_6')
// (17, 6, 'sp4_v_t_44')
// (17, 7, 'sp4_v_b_44')
// (17, 8, 'sp4_v_b_33')
// (17, 9, 'local_g1_4')
// (17, 9, 'lutff_4/in_3')
// (17, 9, 'sp4_v_b_20')
// (17, 10, 'sp4_v_b_9')
// (17, 10, 'sp4_v_t_43')
// (17, 11, 'sp4_v_b_43')
// (17, 12, 'sp4_v_b_30')
// (17, 13, 'neigh_op_tnr_6')
// (17, 13, 'sp4_v_b_19')
// (17, 14, 'neigh_op_rgt_6')
// (17, 14, 'sp4_h_r_1')
// (17, 14, 'sp4_v_b_6')
// (17, 15, 'neigh_op_bnr_6')
// (18, 13, 'neigh_op_top_6')
// (18, 14, 'lutff_6/out')
// (18, 14, 'sp4_h_r_12')
// (18, 15, 'neigh_op_bot_6')
// (19, 13, 'neigh_op_tnl_6')
// (19, 14, 'neigh_op_lft_6')
// (19, 14, 'sp4_h_r_25')
// (19, 15, 'neigh_op_bnl_6')
// (20, 14, 'sp4_h_r_36')
// (21, 14, 'sp4_h_l_36')

reg n1054 = 0;
// (16, 9, 'sp4_r_v_b_44')
// (16, 10, 'local_g0_2')
// (16, 10, 'lutff_3/in_3')
// (16, 10, 'sp4_r_v_b_33')
// (16, 11, 'sp4_r_v_b_20')
// (16, 12, 'sp4_r_v_b_9')
// (17, 8, 'sp4_v_t_44')
// (17, 9, 'sp4_v_b_44')
// (17, 10, 'sp4_v_b_33')
// (17, 11, 'sp4_v_b_20')
// (17, 12, 'sp4_h_r_4')
// (17, 12, 'sp4_v_b_9')
// (18, 12, 'sp4_h_r_17')
// (19, 12, 'sp4_h_r_28')
// (20, 12, 'sp4_h_r_41')
// (20, 13, 'sp4_r_v_b_41')
// (20, 14, 'sp4_r_v_b_28')
// (20, 15, 'sp4_r_v_b_17')
// (20, 16, 'sp4_r_v_b_4')
// (20, 17, 'sp4_r_v_b_36')
// (20, 18, 'neigh_op_tnr_6')
// (20, 18, 'sp4_r_v_b_25')
// (20, 19, 'neigh_op_rgt_6')
// (20, 19, 'sp4_r_v_b_12')
// (20, 20, 'neigh_op_bnr_6')
// (20, 20, 'sp4_r_v_b_1')
// (21, 12, 'sp4_h_l_41')
// (21, 12, 'sp4_v_t_41')
// (21, 13, 'sp4_v_b_41')
// (21, 14, 'sp4_v_b_28')
// (21, 15, 'sp4_v_b_17')
// (21, 16, 'sp4_v_b_4')
// (21, 16, 'sp4_v_t_36')
// (21, 17, 'sp4_v_b_36')
// (21, 18, 'neigh_op_top_6')
// (21, 18, 'sp4_v_b_25')
// (21, 19, 'lutff_6/out')
// (21, 19, 'sp4_v_b_12')
// (21, 20, 'neigh_op_bot_6')
// (21, 20, 'sp4_v_b_1')
// (22, 18, 'neigh_op_tnl_6')
// (22, 19, 'neigh_op_lft_6')
// (22, 20, 'neigh_op_bnl_6')

reg n1055 = 0;
// (16, 10, 'local_g1_2')
// (16, 10, 'lutff_2/in_3')
// (16, 10, 'sp4_h_r_10')
// (17, 10, 'sp4_h_r_23')
// (18, 10, 'sp4_h_r_34')
// (19, 10, 'sp4_h_r_47')
// (19, 11, 'sp4_r_v_b_41')
// (19, 12, 'sp4_r_v_b_28')
// (19, 13, 'neigh_op_tnr_2')
// (19, 13, 'sp4_r_v_b_17')
// (19, 14, 'neigh_op_rgt_2')
// (19, 14, 'sp4_r_v_b_4')
// (19, 15, 'neigh_op_bnr_2')
// (20, 10, 'sp4_h_l_47')
// (20, 10, 'sp4_v_t_41')
// (20, 11, 'sp4_v_b_41')
// (20, 12, 'sp4_v_b_28')
// (20, 13, 'neigh_op_top_2')
// (20, 13, 'sp4_v_b_17')
// (20, 14, 'lutff_2/out')
// (20, 14, 'sp4_v_b_4')
// (20, 15, 'neigh_op_bot_2')
// (21, 13, 'neigh_op_tnl_2')
// (21, 14, 'neigh_op_lft_2')
// (21, 15, 'neigh_op_bnl_2')

reg n1056 = 0;
// (16, 10, 'local_g3_2')
// (16, 10, 'lutff_4/in_3')
// (16, 10, 'sp4_r_v_b_42')
// (16, 11, 'sp4_r_v_b_31')
// (16, 12, 'sp4_r_v_b_18')
// (16, 13, 'sp4_r_v_b_7')
// (17, 9, 'sp4_v_t_42')
// (17, 10, 'sp4_v_b_42')
// (17, 11, 'sp4_v_b_31')
// (17, 12, 'sp4_v_b_18')
// (17, 13, 'sp4_h_r_7')
// (17, 13, 'sp4_v_b_7')
// (18, 13, 'sp4_h_r_18')
// (19, 13, 'sp4_h_r_31')
// (20, 13, 'sp4_h_r_42')
// (20, 14, 'sp4_r_v_b_42')
// (20, 15, 'sp4_r_v_b_31')
// (20, 16, 'sp4_r_v_b_18')
// (20, 17, 'sp4_r_v_b_7')
// (21, 13, 'sp4_h_l_42')
// (21, 13, 'sp4_v_t_42')
// (21, 14, 'sp4_v_b_42')
// (21, 15, 'sp4_v_b_31')
// (21, 16, 'neigh_op_tnr_1')
// (21, 16, 'sp4_v_b_18')
// (21, 17, 'neigh_op_rgt_1')
// (21, 17, 'sp4_h_r_7')
// (21, 17, 'sp4_v_b_7')
// (21, 18, 'neigh_op_bnr_1')
// (22, 16, 'neigh_op_top_1')
// (22, 17, 'lutff_1/out')
// (22, 17, 'sp4_h_r_18')
// (22, 18, 'neigh_op_bot_1')
// (23, 16, 'neigh_op_tnl_1')
// (23, 17, 'neigh_op_lft_1')
// (23, 17, 'sp4_h_r_31')
// (23, 18, 'neigh_op_bnl_1')
// (24, 17, 'sp4_h_r_42')
// (25, 17, 'sp4_h_l_42')

wire n1057;
// (16, 10, 'neigh_op_tnr_0')
// (16, 11, 'neigh_op_rgt_0')
// (16, 12, 'neigh_op_bnr_0')
// (17, 10, 'neigh_op_top_0')
// (17, 11, 'local_g1_0')
// (17, 11, 'lutff_0/out')
// (17, 11, 'lutff_2/in_3')
// (17, 12, 'neigh_op_bot_0')
// (18, 10, 'neigh_op_tnl_0')
// (18, 11, 'neigh_op_lft_0')
// (18, 12, 'neigh_op_bnl_0')

wire n1058;
// (16, 10, 'neigh_op_tnr_2')
// (16, 11, 'neigh_op_rgt_2')
// (16, 11, 'sp4_r_v_b_36')
// (16, 12, 'neigh_op_bnr_2')
// (16, 12, 'sp4_r_v_b_25')
// (16, 13, 'sp4_r_v_b_12')
// (16, 14, 'sp4_r_v_b_1')
// (16, 15, 'sp4_r_v_b_36')
// (16, 16, 'sp4_r_v_b_25')
// (16, 17, 'sp4_r_v_b_12')
// (16, 18, 'sp4_r_v_b_1')
// (17, 10, 'neigh_op_top_2')
// (17, 10, 'sp4_v_t_36')
// (17, 11, 'lutff_2/out')
// (17, 11, 'sp4_v_b_36')
// (17, 12, 'neigh_op_bot_2')
// (17, 12, 'sp4_v_b_25')
// (17, 13, 'sp4_v_b_12')
// (17, 14, 'sp4_v_b_1')
// (17, 14, 'sp4_v_t_36')
// (17, 15, 'sp4_v_b_36')
// (17, 16, 'sp4_v_b_25')
// (17, 17, 'sp4_v_b_12')
// (17, 18, 'sp4_h_r_7')
// (17, 18, 'sp4_v_b_1')
// (18, 10, 'neigh_op_tnl_2')
// (18, 11, 'neigh_op_lft_2')
// (18, 12, 'neigh_op_bnl_2')
// (18, 18, 'sp4_h_r_18')
// (19, 18, 'local_g3_7')
// (19, 18, 'lutff_5/in_1')
// (19, 18, 'sp4_h_r_31')
// (20, 18, 'sp4_h_r_42')
// (21, 18, 'sp4_h_l_42')

wire n1059;
// (16, 10, 'neigh_op_tnr_4')
// (16, 11, 'neigh_op_rgt_4')
// (16, 11, 'sp4_r_v_b_40')
// (16, 12, 'neigh_op_bnr_4')
// (16, 12, 'sp4_r_v_b_29')
// (16, 13, 'sp4_r_v_b_16')
// (16, 14, 'sp4_r_v_b_5')
// (17, 10, 'neigh_op_top_4')
// (17, 10, 'sp4_v_t_40')
// (17, 11, 'lutff_4/out')
// (17, 11, 'sp4_v_b_40')
// (17, 12, 'neigh_op_bot_4')
// (17, 12, 'sp4_v_b_29')
// (17, 13, 'sp4_v_b_16')
// (17, 14, 'sp4_h_r_11')
// (17, 14, 'sp4_v_b_5')
// (18, 10, 'neigh_op_tnl_4')
// (18, 11, 'neigh_op_lft_4')
// (18, 12, 'neigh_op_bnl_4')
// (18, 14, 'sp4_h_r_22')
// (19, 14, 'local_g3_3')
// (19, 14, 'lutff_5/in_1')
// (19, 14, 'sp4_h_r_35')
// (20, 14, 'sp4_h_r_46')
// (21, 14, 'sp4_h_l_46')

wire n1060;
// (16, 10, 'neigh_op_tnr_5')
// (16, 11, 'neigh_op_rgt_5')
// (16, 12, 'neigh_op_bnr_5')
// (17, 10, 'neigh_op_top_5')
// (17, 11, 'local_g2_5')
// (17, 11, 'lutff_4/in_3')
// (17, 11, 'lutff_5/out')
// (17, 12, 'neigh_op_bot_5')
// (18, 10, 'neigh_op_tnl_5')
// (18, 11, 'neigh_op_lft_5')
// (18, 12, 'neigh_op_bnl_5')

reg n1061 = 0;
// (16, 10, 'neigh_op_tnr_6')
// (16, 11, 'neigh_op_rgt_6')
// (16, 12, 'neigh_op_bnr_6')
// (17, 10, 'neigh_op_top_6')
// (17, 11, 'local_g2_6')
// (17, 11, 'lutff_1/in_3')
// (17, 11, 'lutff_6/out')
// (17, 12, 'neigh_op_bot_6')
// (18, 10, 'neigh_op_tnl_6')
// (18, 11, 'neigh_op_lft_6')
// (18, 12, 'neigh_op_bnl_6')

reg n1062 = 0;
// (16, 10, 'neigh_op_tnr_7')
// (16, 11, 'neigh_op_rgt_7')
// (16, 12, 'neigh_op_bnr_7')
// (17, 10, 'neigh_op_top_7')
// (17, 11, 'local_g1_7')
// (17, 11, 'lutff_3/in_3')
// (17, 11, 'lutff_7/out')
// (17, 12, 'neigh_op_bot_7')
// (18, 10, 'neigh_op_tnl_7')
// (18, 11, 'neigh_op_lft_7')
// (18, 12, 'neigh_op_bnl_7')

reg n1063 = 0;
// (16, 11, 'neigh_op_tnr_0')
// (16, 12, 'neigh_op_rgt_0')
// (16, 13, 'neigh_op_bnr_0')
// (17, 11, 'neigh_op_top_0')
// (17, 12, 'local_g1_0')
// (17, 12, 'lutff_0/out')
// (17, 12, 'lutff_2/in_3')
// (17, 13, 'neigh_op_bot_0')
// (18, 11, 'neigh_op_tnl_0')
// (18, 12, 'neigh_op_lft_0')
// (18, 13, 'neigh_op_bnl_0')

wire n1064;
// (16, 11, 'neigh_op_tnr_2')
// (16, 12, 'neigh_op_rgt_2')
// (16, 13, 'neigh_op_bnr_2')
// (17, 11, 'neigh_op_top_2')
// (17, 12, 'lutff_2/out')
// (17, 13, 'neigh_op_bot_2')
// (18, 11, 'neigh_op_tnl_2')
// (18, 12, 'neigh_op_lft_2')
// (18, 13, 'local_g3_2')
// (18, 13, 'lutff_6/in_3')
// (18, 13, 'neigh_op_bnl_2')

wire n1065;
// (16, 11, 'neigh_op_tnr_3')
// (16, 12, 'neigh_op_rgt_3')
// (16, 13, 'neigh_op_bnr_3')
// (17, 11, 'neigh_op_top_3')
// (17, 12, 'lutff_3/out')
// (17, 13, 'local_g1_3')
// (17, 13, 'lutff_3/in_3')
// (17, 13, 'neigh_op_bot_3')
// (18, 11, 'neigh_op_tnl_3')
// (18, 12, 'neigh_op_lft_3')
// (18, 13, 'neigh_op_bnl_3')

wire n1066;
// (16, 11, 'neigh_op_tnr_4')
// (16, 12, 'neigh_op_rgt_4')
// (16, 13, 'neigh_op_bnr_4')
// (17, 11, 'neigh_op_top_4')
// (17, 12, 'lutff_4/out')
// (17, 13, 'local_g0_4')
// (17, 13, 'lutff_3/in_1')
// (17, 13, 'neigh_op_bot_4')
// (18, 11, 'neigh_op_tnl_4')
// (18, 12, 'neigh_op_lft_4')
// (18, 13, 'neigh_op_bnl_4')

wire n1067;
// (16, 11, 'neigh_op_tnr_5')
// (16, 12, 'neigh_op_rgt_5')
// (16, 13, 'neigh_op_bnr_5')
// (17, 11, 'neigh_op_top_5')
// (17, 12, 'lutff_5/out')
// (17, 12, 'sp4_r_v_b_43')
// (17, 13, 'neigh_op_bot_5')
// (17, 13, 'sp4_r_v_b_30')
// (17, 14, 'sp4_r_v_b_19')
// (17, 15, 'sp4_r_v_b_6')
// (18, 11, 'neigh_op_tnl_5')
// (18, 11, 'sp4_v_t_43')
// (18, 12, 'neigh_op_lft_5')
// (18, 12, 'sp4_v_b_43')
// (18, 13, 'neigh_op_bnl_5')
// (18, 13, 'sp4_v_b_30')
// (18, 14, 'local_g0_3')
// (18, 14, 'lutff_5/in_0')
// (18, 14, 'sp4_v_b_19')
// (18, 15, 'sp4_v_b_6')

wire n1068;
// (16, 11, 'neigh_op_tnr_6')
// (16, 11, 'sp4_r_v_b_41')
// (16, 12, 'neigh_op_rgt_6')
// (16, 12, 'sp4_r_v_b_28')
// (16, 13, 'neigh_op_bnr_6')
// (16, 13, 'sp4_r_v_b_17')
// (16, 14, 'sp4_r_v_b_4')
// (17, 10, 'sp4_v_t_41')
// (17, 11, 'neigh_op_top_6')
// (17, 11, 'sp4_v_b_41')
// (17, 12, 'lutff_6/out')
// (17, 12, 'sp4_v_b_28')
// (17, 13, 'neigh_op_bot_6')
// (17, 13, 'sp4_v_b_17')
// (17, 14, 'sp4_h_r_4')
// (17, 14, 'sp4_v_b_4')
// (18, 11, 'neigh_op_tnl_6')
// (18, 12, 'neigh_op_lft_6')
// (18, 13, 'neigh_op_bnl_6')
// (18, 14, 'sp4_h_r_17')
// (19, 14, 'sp4_h_r_28')
// (20, 14, 'local_g2_1')
// (20, 14, 'lutff_4/in_3')
// (20, 14, 'sp4_h_r_41')
// (21, 14, 'sp4_h_l_41')

wire n1069;
// (16, 11, 'neigh_op_tnr_7')
// (16, 12, 'neigh_op_rgt_7')
// (16, 12, 'sp4_r_v_b_46')
// (16, 13, 'neigh_op_bnr_7')
// (16, 13, 'sp4_r_v_b_35')
// (16, 14, 'sp4_r_v_b_22')
// (16, 15, 'sp4_r_v_b_11')
// (17, 11, 'neigh_op_top_7')
// (17, 11, 'sp4_v_t_46')
// (17, 12, 'lutff_7/out')
// (17, 12, 'sp4_v_b_46')
// (17, 13, 'neigh_op_bot_7')
// (17, 13, 'sp4_v_b_35')
// (17, 14, 'sp4_v_b_22')
// (17, 15, 'sp4_h_r_5')
// (17, 15, 'sp4_v_b_11')
// (18, 11, 'neigh_op_tnl_7')
// (18, 12, 'neigh_op_lft_7')
// (18, 13, 'neigh_op_bnl_7')
// (18, 15, 'sp4_h_r_16')
// (19, 15, 'sp4_h_r_29')
// (20, 15, 'sp4_h_r_40')
// (20, 16, 'sp4_r_v_b_40')
// (20, 17, 'sp4_r_v_b_29')
// (20, 18, 'sp4_r_v_b_16')
// (20, 19, 'sp4_r_v_b_5')
// (21, 15, 'sp4_h_l_40')
// (21, 15, 'sp4_v_t_40')
// (21, 16, 'sp4_v_b_40')
// (21, 17, 'sp4_v_b_29')
// (21, 18, 'sp4_v_b_16')
// (21, 19, 'local_g1_5')
// (21, 19, 'lutff_1/in_3')
// (21, 19, 'sp4_v_b_5')

wire n1070;
// (16, 12, 'lutff_2/lout')
// (16, 12, 'lutff_3/in_2')

wire n1071;
// (16, 12, 'lutff_3/lout')
// (16, 12, 'lutff_4/in_2')

wire n1072;
// (16, 12, 'lutff_6/lout')
// (16, 12, 'lutff_7/in_2')

reg n1073 = 0;
// (16, 12, 'neigh_op_tnr_0')
// (16, 13, 'neigh_op_rgt_0')
// (16, 14, 'neigh_op_bnr_0')
// (17, 12, 'neigh_op_top_0')
// (17, 13, 'local_g1_0')
// (17, 13, 'lutff_0/out')
// (17, 13, 'lutff_2/in_3')
// (17, 14, 'neigh_op_bot_0')
// (18, 12, 'neigh_op_tnl_0')
// (18, 13, 'neigh_op_lft_0')
// (18, 14, 'neigh_op_bnl_0')

wire n1074;
// (16, 12, 'neigh_op_tnr_2')
// (16, 13, 'neigh_op_rgt_2')
// (16, 14, 'neigh_op_bnr_2')
// (17, 12, 'neigh_op_top_2')
// (17, 13, 'lutff_2/out')
// (17, 14, 'neigh_op_bot_2')
// (18, 12, 'neigh_op_tnl_2')
// (18, 13, 'local_g1_2')
// (18, 13, 'lutff_6/in_1')
// (18, 13, 'neigh_op_lft_2')
// (18, 14, 'neigh_op_bnl_2')

wire n1075;
// (16, 12, 'neigh_op_tnr_5')
// (16, 13, 'neigh_op_rgt_5')
// (16, 13, 'sp4_r_v_b_42')
// (16, 14, 'neigh_op_bnr_5')
// (16, 14, 'sp4_r_v_b_31')
// (16, 15, 'sp4_r_v_b_18')
// (16, 16, 'sp4_r_v_b_7')
// (17, 12, 'neigh_op_top_5')
// (17, 12, 'sp4_v_t_42')
// (17, 13, 'lutff_5/out')
// (17, 13, 'sp4_v_b_42')
// (17, 14, 'neigh_op_bot_5')
// (17, 14, 'sp4_v_b_31')
// (17, 15, 'sp4_v_b_18')
// (17, 16, 'local_g0_7')
// (17, 16, 'lutff_4/in_3')
// (17, 16, 'sp4_v_b_7')
// (18, 12, 'neigh_op_tnl_5')
// (18, 13, 'neigh_op_lft_5')
// (18, 14, 'neigh_op_bnl_5')

wire n1076;
// (16, 12, 'neigh_op_tnr_7')
// (16, 13, 'neigh_op_rgt_7')
// (16, 14, 'neigh_op_bnr_7')
// (17, 12, 'neigh_op_top_7')
// (17, 13, 'local_g2_7')
// (17, 13, 'lutff_4/in_1')
// (17, 13, 'lutff_7/out')
// (17, 14, 'neigh_op_bot_7')
// (18, 12, 'neigh_op_tnl_7')
// (18, 13, 'neigh_op_lft_7')
// (18, 14, 'neigh_op_bnl_7')

wire n1077;
// (16, 12, 'sp4_h_r_7')
// (17, 12, 'sp4_h_r_18')
// (18, 11, 'neigh_op_tnr_5')
// (18, 12, 'neigh_op_rgt_5')
// (18, 12, 'sp4_h_r_31')
// (18, 13, 'neigh_op_bnr_5')
// (19, 11, 'neigh_op_top_5')
// (19, 12, 'lutff_5/out')
// (19, 12, 'sp4_h_r_42')
// (19, 13, 'neigh_op_bot_5')
// (20, 11, 'neigh_op_tnl_5')
// (20, 12, 'neigh_op_lft_5')
// (20, 12, 'sp4_h_l_42')
// (20, 12, 'sp4_h_r_10')
// (20, 13, 'neigh_op_bnl_5')
// (21, 12, 'sp4_h_r_23')
// (22, 12, 'local_g2_2')
// (22, 12, 'lutff_global/cen')
// (22, 12, 'sp4_h_r_34')
// (23, 12, 'sp4_h_r_47')
// (24, 12, 'sp4_h_l_47')

reg n1078 = 0;
// (16, 12, 'sp4_r_v_b_39')
// (16, 13, 'sp4_r_v_b_26')
// (16, 14, 'sp4_r_v_b_15')
// (16, 15, 'sp4_r_v_b_2')
// (16, 16, 'sp4_r_v_b_39')
// (16, 17, 'sp4_r_v_b_26')
// (16, 18, 'sp4_r_v_b_15')
// (16, 19, 'sp4_r_v_b_2')
// (17, 11, 'sp4_v_t_39')
// (17, 12, 'sp4_v_b_39')
// (17, 13, 'sp4_v_b_26')
// (17, 14, 'local_g0_7')
// (17, 14, 'lutff_4/in_3')
// (17, 14, 'sp4_v_b_15')
// (17, 15, 'sp4_v_b_2')
// (17, 15, 'sp4_v_t_39')
// (17, 16, 'sp4_v_b_39')
// (17, 17, 'sp4_v_b_26')
// (17, 18, 'sp4_v_b_15')
// (17, 19, 'sp4_h_r_2')
// (17, 19, 'sp4_v_b_2')
// (18, 18, 'neigh_op_tnr_5')
// (18, 19, 'neigh_op_rgt_5')
// (18, 19, 'sp4_h_r_15')
// (18, 20, 'neigh_op_bnr_5')
// (19, 18, 'neigh_op_top_5')
// (19, 19, 'lutff_5/out')
// (19, 19, 'sp4_h_r_26')
// (19, 20, 'neigh_op_bot_5')
// (20, 18, 'neigh_op_tnl_5')
// (20, 19, 'neigh_op_lft_5')
// (20, 19, 'sp4_h_r_39')
// (20, 20, 'neigh_op_bnl_5')
// (21, 19, 'sp4_h_l_39')

wire n1079;
// (16, 13, 'lutff_6/lout')
// (16, 13, 'lutff_7/in_2')

reg n1080 = 0;
// (16, 13, 'neigh_op_tnr_2')
// (16, 14, 'neigh_op_rgt_2')
// (16, 15, 'neigh_op_bnr_2')
// (17, 13, 'neigh_op_top_2')
// (17, 14, 'local_g3_2')
// (17, 14, 'lutff_0/in_3')
// (17, 14, 'lutff_2/out')
// (17, 15, 'neigh_op_bot_2')
// (18, 13, 'neigh_op_tnl_2')
// (18, 14, 'neigh_op_lft_2')
// (18, 15, 'neigh_op_bnl_2')

wire n1081;
// (16, 13, 'neigh_op_tnr_4')
// (16, 14, 'neigh_op_rgt_4')
// (16, 15, 'neigh_op_bnr_4')
// (17, 13, 'neigh_op_top_4')
// (17, 14, 'lutff_4/out')
// (17, 15, 'neigh_op_bot_4')
// (18, 13, 'local_g2_4')
// (18, 13, 'lutff_7/in_1')
// (18, 13, 'neigh_op_tnl_4')
// (18, 14, 'neigh_op_lft_4')
// (18, 15, 'neigh_op_bnl_4')

reg n1082 = 0;
// (16, 13, 'neigh_op_tnr_5')
// (16, 14, 'neigh_op_rgt_5')
// (16, 15, 'neigh_op_bnr_5')
// (17, 13, 'neigh_op_top_5')
// (17, 14, 'local_g1_5')
// (17, 14, 'lutff_3/in_3')
// (17, 14, 'lutff_5/out')
// (17, 15, 'neigh_op_bot_5')
// (18, 13, 'neigh_op_tnl_5')
// (18, 14, 'neigh_op_lft_5')
// (18, 15, 'neigh_op_bnl_5')

wire n1083;
// (16, 13, 'neigh_op_tnr_7')
// (16, 14, 'neigh_op_rgt_7')
// (16, 15, 'neigh_op_bnr_7')
// (17, 13, 'local_g0_7')
// (17, 13, 'lutff_4/in_3')
// (17, 13, 'neigh_op_top_7')
// (17, 14, 'lutff_7/out')
// (17, 15, 'neigh_op_bot_7')
// (18, 13, 'neigh_op_tnl_7')
// (18, 14, 'neigh_op_lft_7')
// (18, 15, 'neigh_op_bnl_7')

wire n1084;
// (16, 13, 'sp4_h_r_0')
// (17, 13, 'sp4_h_r_13')
// (18, 13, 'local_g2_0')
// (18, 13, 'lutff_3/in_3')
// (18, 13, 'sp4_h_r_24')
// (19, 13, 'sp4_h_r_37')
// (19, 14, 'sp4_r_v_b_43')
// (19, 15, 'sp4_r_v_b_30')
// (19, 16, 'sp4_r_v_b_19')
// (19, 17, 'sp4_r_v_b_6')
// (20, 13, 'sp4_h_l_37')
// (20, 13, 'sp4_v_t_43')
// (20, 14, 'sp4_v_b_43')
// (20, 15, 'sp4_v_b_30')
// (20, 16, 'neigh_op_tnr_6')
// (20, 16, 'sp4_v_b_19')
// (20, 17, 'neigh_op_rgt_6')
// (20, 17, 'sp4_h_r_1')
// (20, 17, 'sp4_v_b_6')
// (20, 18, 'neigh_op_bnr_6')
// (21, 16, 'neigh_op_top_6')
// (21, 17, 'lutff_6/out')
// (21, 17, 'sp4_h_r_12')
// (21, 18, 'neigh_op_bot_6')
// (22, 16, 'neigh_op_tnl_6')
// (22, 17, 'neigh_op_lft_6')
// (22, 17, 'sp4_h_r_25')
// (22, 18, 'neigh_op_bnl_6')
// (23, 17, 'sp4_h_r_36')
// (24, 17, 'sp4_h_l_36')

reg n1085 = 0;
// (16, 13, 'sp4_h_r_7')
// (17, 13, 'local_g1_2')
// (17, 13, 'lutff_2/in_1')
// (17, 13, 'sp4_h_r_18')
// (18, 13, 'sp4_h_r_31')
// (19, 13, 'sp4_h_r_42')
// (19, 14, 'sp4_r_v_b_36')
// (19, 15, 'neigh_op_tnr_6')
// (19, 15, 'sp4_r_v_b_25')
// (19, 16, 'neigh_op_rgt_6')
// (19, 16, 'sp4_r_v_b_12')
// (19, 17, 'neigh_op_bnr_6')
// (19, 17, 'sp4_r_v_b_1')
// (20, 13, 'sp4_h_l_42')
// (20, 13, 'sp4_v_t_36')
// (20, 14, 'sp4_v_b_36')
// (20, 15, 'neigh_op_top_6')
// (20, 15, 'sp4_v_b_25')
// (20, 16, 'lutff_6/out')
// (20, 16, 'sp4_v_b_12')
// (20, 17, 'neigh_op_bot_6')
// (20, 17, 'sp4_v_b_1')
// (21, 15, 'neigh_op_tnl_6')
// (21, 16, 'neigh_op_lft_6')
// (21, 17, 'neigh_op_bnl_6')

wire n1086;
// (16, 14, 'lutff_5/lout')
// (16, 14, 'lutff_6/in_2')

wire n1087;
// (16, 14, 'neigh_op_tnr_1')
// (16, 15, 'neigh_op_rgt_1')
// (16, 16, 'neigh_op_bnr_1')
// (17, 12, 'sp4_r_v_b_38')
// (17, 13, 'sp4_r_v_b_27')
// (17, 14, 'neigh_op_top_1')
// (17, 14, 'sp4_r_v_b_14')
// (17, 15, 'lutff_1/out')
// (17, 15, 'sp4_r_v_b_3')
// (17, 16, 'neigh_op_bot_1')
// (18, 11, 'sp4_v_t_38')
// (18, 12, 'sp4_v_b_38')
// (18, 13, 'local_g3_3')
// (18, 13, 'lutff_7/in_3')
// (18, 13, 'sp4_v_b_27')
// (18, 14, 'neigh_op_tnl_1')
// (18, 14, 'sp4_v_b_14')
// (18, 15, 'neigh_op_lft_1')
// (18, 15, 'sp4_v_b_3')
// (18, 16, 'neigh_op_bnl_1')

reg n1088 = 0;
// (16, 14, 'neigh_op_tnr_2')
// (16, 15, 'neigh_op_rgt_2')
// (16, 16, 'neigh_op_bnr_2')
// (17, 14, 'neigh_op_top_2')
// (17, 15, 'local_g3_2')
// (17, 15, 'lutff_0/in_3')
// (17, 15, 'lutff_2/out')
// (17, 16, 'neigh_op_bot_2')
// (18, 14, 'neigh_op_tnl_2')
// (18, 15, 'neigh_op_lft_2')
// (18, 16, 'neigh_op_bnl_2')

wire n1089;
// (16, 14, 'neigh_op_tnr_4')
// (16, 15, 'neigh_op_rgt_4')
// (16, 16, 'neigh_op_bnr_4')
// (17, 14, 'neigh_op_top_4')
// (17, 15, 'lutff_4/out')
// (17, 16, 'local_g0_4')
// (17, 16, 'lutff_6/in_0')
// (17, 16, 'neigh_op_bot_4')
// (18, 14, 'neigh_op_tnl_4')
// (18, 15, 'neigh_op_lft_4')
// (18, 16, 'neigh_op_bnl_4')

wire n1090;
// (16, 14, 'neigh_op_tnr_6')
// (16, 15, 'neigh_op_rgt_6')
// (16, 16, 'neigh_op_bnr_6')
// (17, 14, 'neigh_op_top_6')
// (17, 15, 'lutff_6/out')
// (17, 16, 'neigh_op_bot_6')
// (18, 14, 'local_g2_6')
// (18, 14, 'lutff_3/in_1')
// (18, 14, 'neigh_op_tnl_6')
// (18, 15, 'neigh_op_lft_6')
// (18, 16, 'neigh_op_bnl_6')

wire n1091;
// (16, 14, 'neigh_op_tnr_7')
// (16, 15, 'neigh_op_rgt_7')
// (16, 15, 'sp4_r_v_b_46')
// (16, 16, 'neigh_op_bnr_7')
// (16, 16, 'sp4_r_v_b_35')
// (16, 17, 'sp4_r_v_b_22')
// (16, 18, 'sp4_r_v_b_11')
// (17, 14, 'neigh_op_top_7')
// (17, 14, 'sp4_v_t_46')
// (17, 15, 'lutff_7/out')
// (17, 15, 'sp4_v_b_46')
// (17, 16, 'neigh_op_bot_7')
// (17, 16, 'sp4_v_b_35')
// (17, 17, 'local_g1_6')
// (17, 17, 'lutff_0/in_3')
// (17, 17, 'sp4_v_b_22')
// (17, 18, 'sp4_v_b_11')
// (18, 14, 'neigh_op_tnl_7')
// (18, 15, 'neigh_op_lft_7')
// (18, 16, 'neigh_op_bnl_7')

wire n1092;
// (16, 14, 'sp12_h_r_1')
// (17, 14, 'sp12_h_r_2')
// (18, 14, 'local_g1_5')
// (18, 14, 'lutff_3/in_3')
// (18, 14, 'sp12_h_r_5')
// (19, 14, 'sp12_h_r_6')
// (20, 13, 'neigh_op_tnr_1')
// (20, 14, 'neigh_op_rgt_1')
// (20, 14, 'sp12_h_r_9')
// (20, 15, 'neigh_op_bnr_1')
// (21, 13, 'neigh_op_top_1')
// (21, 14, 'lutff_1/out')
// (21, 14, 'sp12_h_r_10')
// (21, 15, 'neigh_op_bot_1')
// (22, 13, 'neigh_op_tnl_1')
// (22, 14, 'neigh_op_lft_1')
// (22, 14, 'sp12_h_r_13')
// (22, 15, 'neigh_op_bnl_1')
// (23, 14, 'sp12_h_r_14')
// (24, 14, 'sp12_h_r_17')
// (25, 14, 'sp12_h_r_18')
// (26, 14, 'sp12_h_r_21')
// (27, 14, 'sp12_h_r_22')
// (28, 14, 'sp12_h_l_22')

wire n1093;
// (16, 14, 'sp4_h_r_0')
// (17, 14, 'sp4_h_r_13')
// (18, 14, 'local_g2_0')
// (18, 14, 'lutff_5/in_3')
// (18, 14, 'sp4_h_r_24')
// (19, 14, 'sp4_h_r_37')
// (19, 15, 'sp4_r_v_b_37')
// (19, 16, 'sp4_r_v_b_24')
// (19, 17, 'neigh_op_tnr_0')
// (19, 17, 'sp4_r_v_b_13')
// (19, 18, 'neigh_op_rgt_0')
// (19, 18, 'sp4_r_v_b_0')
// (19, 19, 'neigh_op_bnr_0')
// (20, 14, 'sp4_h_l_37')
// (20, 14, 'sp4_v_t_37')
// (20, 15, 'sp4_v_b_37')
// (20, 16, 'sp4_v_b_24')
// (20, 17, 'neigh_op_top_0')
// (20, 17, 'sp4_v_b_13')
// (20, 18, 'lutff_0/out')
// (20, 18, 'sp4_v_b_0')
// (20, 19, 'neigh_op_bot_0')
// (21, 17, 'neigh_op_tnl_0')
// (21, 18, 'neigh_op_lft_0')
// (21, 19, 'neigh_op_bnl_0')

wire n1094;
// (16, 14, 'sp4_h_r_11')
// (17, 14, 'sp4_h_r_22')
// (18, 14, 'local_g2_3')
// (18, 14, 'lutff_4/in_3')
// (18, 14, 'sp4_h_r_35')
// (19, 14, 'sp4_h_r_46')
// (19, 15, 'sp4_r_v_b_40')
// (19, 16, 'neigh_op_tnr_0')
// (19, 16, 'sp4_r_v_b_29')
// (19, 17, 'neigh_op_rgt_0')
// (19, 17, 'sp4_r_v_b_16')
// (19, 18, 'neigh_op_bnr_0')
// (19, 18, 'sp4_r_v_b_5')
// (20, 14, 'sp4_h_l_46')
// (20, 14, 'sp4_v_t_40')
// (20, 15, 'sp4_v_b_40')
// (20, 16, 'neigh_op_top_0')
// (20, 16, 'sp4_v_b_29')
// (20, 17, 'lutff_0/out')
// (20, 17, 'sp4_v_b_16')
// (20, 18, 'neigh_op_bot_0')
// (20, 18, 'sp4_v_b_5')
// (21, 16, 'neigh_op_tnl_0')
// (21, 17, 'neigh_op_lft_0')
// (21, 18, 'neigh_op_bnl_0')

reg n1095 = 0;
// (16, 14, 'sp4_h_r_7')
// (17, 14, 'sp4_h_r_18')
// (18, 14, 'sp4_h_r_31')
// (19, 10, 'neigh_op_tnr_5')
// (19, 11, 'neigh_op_rgt_5')
// (19, 11, 'sp4_r_v_b_42')
// (19, 12, 'neigh_op_bnr_5')
// (19, 12, 'sp4_r_v_b_31')
// (19, 13, 'sp4_r_v_b_18')
// (19, 14, 'local_g3_2')
// (19, 14, 'lutff_3/in_0')
// (19, 14, 'sp4_h_r_42')
// (19, 14, 'sp4_r_v_b_7')
// (20, 10, 'neigh_op_top_5')
// (20, 10, 'sp4_v_t_42')
// (20, 11, 'lutff_5/out')
// (20, 11, 'sp4_v_b_42')
// (20, 12, 'neigh_op_bot_5')
// (20, 12, 'sp4_v_b_31')
// (20, 13, 'sp4_v_b_18')
// (20, 14, 'sp4_h_l_42')
// (20, 14, 'sp4_v_b_7')
// (21, 10, 'neigh_op_tnl_5')
// (21, 11, 'neigh_op_lft_5')
// (21, 12, 'neigh_op_bnl_5')

reg n1096 = 0;
// (16, 14, 'sp4_h_r_9')
// (17, 14, 'local_g1_4')
// (17, 14, 'lutff_6/in_3')
// (17, 14, 'sp4_h_r_20')
// (18, 14, 'sp4_h_r_33')
// (19, 10, 'neigh_op_tnr_6')
// (19, 11, 'neigh_op_rgt_6')
// (19, 11, 'sp4_r_v_b_44')
// (19, 12, 'neigh_op_bnr_6')
// (19, 12, 'sp4_r_v_b_33')
// (19, 13, 'sp4_r_v_b_20')
// (19, 14, 'sp4_h_r_44')
// (19, 14, 'sp4_r_v_b_9')
// (20, 10, 'neigh_op_top_6')
// (20, 10, 'sp4_v_t_44')
// (20, 11, 'lutff_6/out')
// (20, 11, 'sp4_v_b_44')
// (20, 12, 'neigh_op_bot_6')
// (20, 12, 'sp4_v_b_33')
// (20, 13, 'sp4_v_b_20')
// (20, 14, 'sp4_h_l_44')
// (20, 14, 'sp4_v_b_9')
// (21, 10, 'neigh_op_tnl_6')
// (21, 11, 'neigh_op_lft_6')
// (21, 12, 'neigh_op_bnl_6')

wire n1097;
// (16, 15, 'lutff_0/lout')
// (16, 15, 'lutff_1/in_2')

wire n1098;
// (16, 15, 'lutff_3/lout')
// (16, 15, 'lutff_4/in_2')

wire n1099;
// (16, 15, 'lutff_6/lout')
// (16, 15, 'lutff_7/in_2')

wire n1100;
// (16, 15, 'neigh_op_tnr_0')
// (16, 16, 'neigh_op_rgt_0')
// (16, 17, 'neigh_op_bnr_0')
// (17, 15, 'neigh_op_top_0')
// (17, 16, 'local_g2_0')
// (17, 16, 'lutff_0/out')
// (17, 16, 'lutff_5/in_3')
// (17, 17, 'neigh_op_bot_0')
// (18, 15, 'neigh_op_tnl_0')
// (18, 16, 'neigh_op_lft_0')
// (18, 17, 'neigh_op_bnl_0')

wire n1101;
// (16, 15, 'neigh_op_tnr_1')
// (16, 16, 'neigh_op_rgt_1')
// (16, 17, 'neigh_op_bnr_1')
// (17, 15, 'neigh_op_top_1')
// (17, 16, 'local_g2_1')
// (17, 16, 'lutff_0/in_3')
// (17, 16, 'lutff_1/out')
// (17, 17, 'neigh_op_bot_1')
// (18, 15, 'neigh_op_tnl_1')
// (18, 16, 'neigh_op_lft_1')
// (18, 17, 'neigh_op_bnl_1')

wire n1102;
// (16, 15, 'neigh_op_tnr_3')
// (16, 16, 'neigh_op_rgt_3')
// (16, 17, 'neigh_op_bnr_3')
// (17, 15, 'neigh_op_top_3')
// (17, 16, 'local_g0_3')
// (17, 16, 'lutff_3/out')
// (17, 16, 'lutff_6/in_3')
// (17, 17, 'neigh_op_bot_3')
// (18, 15, 'neigh_op_tnl_3')
// (18, 16, 'neigh_op_lft_3')
// (18, 17, 'neigh_op_bnl_3')

reg n1103 = 0;
// (16, 15, 'sp4_h_r_2')
// (17, 15, 'local_g1_7')
// (17, 15, 'lutff_1/in_3')
// (17, 15, 'sp4_h_r_15')
// (18, 15, 'sp4_h_r_26')
// (19, 11, 'neigh_op_tnr_6')
// (19, 12, 'neigh_op_rgt_6')
// (19, 12, 'sp4_r_v_b_44')
// (19, 13, 'neigh_op_bnr_6')
// (19, 13, 'sp4_r_v_b_33')
// (19, 14, 'sp4_r_v_b_20')
// (19, 15, 'sp4_h_r_39')
// (19, 15, 'sp4_r_v_b_9')
// (20, 11, 'neigh_op_top_6')
// (20, 11, 'sp4_v_t_44')
// (20, 12, 'lutff_6/out')
// (20, 12, 'sp4_v_b_44')
// (20, 13, 'neigh_op_bot_6')
// (20, 13, 'sp4_v_b_33')
// (20, 14, 'sp4_v_b_20')
// (20, 15, 'sp4_h_l_39')
// (20, 15, 'sp4_v_b_9')
// (21, 11, 'neigh_op_tnl_6')
// (21, 12, 'neigh_op_lft_6')
// (21, 13, 'neigh_op_bnl_6')

reg n1104 = 0;
// (16, 15, 'sp4_h_r_8')
// (17, 15, 'sp4_h_r_21')
// (18, 15, 'local_g3_0')
// (18, 15, 'lutff_2/in_3')
// (18, 15, 'sp4_h_r_32')
// (19, 15, 'sp4_h_r_45')
// (20, 15, 'sp4_h_l_45')
// (20, 15, 'sp4_h_r_5')
// (21, 15, 'sp4_h_r_16')
// (22, 15, 'sp4_h_r_29')
// (23, 12, 'sp4_r_v_b_40')
// (23, 13, 'neigh_op_tnr_0')
// (23, 13, 'sp4_r_v_b_29')
// (23, 14, 'neigh_op_rgt_0')
// (23, 14, 'sp4_r_v_b_16')
// (23, 15, 'neigh_op_bnr_0')
// (23, 15, 'sp4_h_r_40')
// (23, 15, 'sp4_r_v_b_5')
// (24, 11, 'sp4_v_t_40')
// (24, 12, 'sp4_v_b_40')
// (24, 13, 'neigh_op_top_0')
// (24, 13, 'sp4_v_b_29')
// (24, 14, 'lutff_0/out')
// (24, 14, 'sp4_v_b_16')
// (24, 15, 'neigh_op_bot_0')
// (24, 15, 'sp4_h_l_40')
// (24, 15, 'sp4_v_b_5')
// (25, 13, 'neigh_op_tnl_0')
// (25, 14, 'neigh_op_lft_0')
// (25, 15, 'neigh_op_bnl_0')

wire n1105;
// (16, 15, 'sp4_r_v_b_40')
// (16, 16, 'neigh_op_tnr_0')
// (16, 16, 'sp4_r_v_b_29')
// (16, 17, 'neigh_op_rgt_0')
// (16, 17, 'sp4_r_v_b_16')
// (16, 18, 'neigh_op_bnr_0')
// (16, 18, 'sp4_r_v_b_5')
// (17, 14, 'sp4_h_r_10')
// (17, 14, 'sp4_v_t_40')
// (17, 15, 'sp4_v_b_40')
// (17, 16, 'neigh_op_top_0')
// (17, 16, 'sp4_v_b_29')
// (17, 17, 'lutff_0/out')
// (17, 17, 'sp4_v_b_16')
// (17, 18, 'neigh_op_bot_0')
// (17, 18, 'sp4_v_b_5')
// (18, 14, 'sp4_h_r_23')
// (18, 16, 'neigh_op_tnl_0')
// (18, 17, 'neigh_op_lft_0')
// (18, 18, 'neigh_op_bnl_0')
// (19, 14, 'sp4_h_r_34')
// (20, 14, 'local_g2_7')
// (20, 14, 'lutff_0/in_1')
// (20, 14, 'sp4_h_r_47')
// (21, 14, 'sp4_h_l_47')

wire n1106;
// (16, 16, 'neigh_op_tnr_2')
// (16, 17, 'neigh_op_rgt_2')
// (16, 18, 'neigh_op_bnr_2')
// (17, 15, 'sp4_r_v_b_45')
// (17, 16, 'neigh_op_top_2')
// (17, 16, 'sp4_r_v_b_32')
// (17, 17, 'lutff_2/out')
// (17, 17, 'sp4_r_v_b_21')
// (17, 18, 'neigh_op_bot_2')
// (17, 18, 'sp4_r_v_b_8')
// (18, 14, 'sp4_v_t_45')
// (18, 15, 'local_g2_5')
// (18, 15, 'lutff_6/in_1')
// (18, 15, 'sp4_v_b_45')
// (18, 16, 'neigh_op_tnl_2')
// (18, 16, 'sp4_v_b_32')
// (18, 17, 'neigh_op_lft_2')
// (18, 17, 'sp4_v_b_21')
// (18, 18, 'neigh_op_bnl_2')
// (18, 18, 'sp4_v_b_8')

wire n1107;
// (16, 16, 'neigh_op_tnr_3')
// (16, 17, 'neigh_op_rgt_3')
// (16, 18, 'neigh_op_bnr_3')
// (17, 16, 'neigh_op_top_3')
// (17, 17, 'local_g0_3')
// (17, 17, 'lutff_2/in_3')
// (17, 17, 'lutff_3/out')
// (17, 18, 'neigh_op_bot_3')
// (18, 16, 'neigh_op_tnl_3')
// (18, 17, 'neigh_op_lft_3')
// (18, 18, 'neigh_op_bnl_3')

reg n1108 = 0;
// (16, 16, 'neigh_op_tnr_4')
// (16, 17, 'neigh_op_rgt_4')
// (16, 18, 'neigh_op_bnr_4')
// (17, 16, 'neigh_op_top_4')
// (17, 17, 'local_g1_4')
// (17, 17, 'lutff_0/in_1')
// (17, 17, 'lutff_4/out')
// (17, 18, 'neigh_op_bot_4')
// (18, 16, 'neigh_op_tnl_4')
// (18, 17, 'neigh_op_lft_4')
// (18, 18, 'neigh_op_bnl_4')

wire n1109;
// (16, 16, 'neigh_op_tnr_6')
// (16, 17, 'neigh_op_rgt_6')
// (16, 17, 'sp4_r_v_b_44')
// (16, 18, 'neigh_op_bnr_6')
// (16, 18, 'sp4_r_v_b_33')
// (16, 19, 'sp4_r_v_b_20')
// (16, 20, 'sp4_r_v_b_9')
// (16, 21, 'sp4_r_v_b_40')
// (16, 22, 'sp4_r_v_b_29')
// (16, 23, 'sp4_r_v_b_16')
// (16, 24, 'sp4_r_v_b_5')
// (16, 25, 'sp4_r_v_b_36')
// (16, 26, 'sp4_r_v_b_25')
// (16, 27, 'sp4_r_v_b_12')
// (16, 28, 'sp4_r_v_b_1')
// (17, 16, 'neigh_op_top_6')
// (17, 16, 'sp4_v_t_44')
// (17, 17, 'lutff_6/out')
// (17, 17, 'sp4_v_b_44')
// (17, 18, 'neigh_op_bot_6')
// (17, 18, 'sp4_v_b_33')
// (17, 19, 'sp4_v_b_20')
// (17, 20, 'sp4_v_b_9')
// (17, 20, 'sp4_v_t_40')
// (17, 21, 'sp4_v_b_40')
// (17, 22, 'sp4_v_b_29')
// (17, 23, 'sp4_v_b_16')
// (17, 24, 'sp4_v_b_5')
// (17, 24, 'sp4_v_t_36')
// (17, 25, 'local_g2_4')
// (17, 25, 'lutff_0/in_0')
// (17, 25, 'sp4_v_b_36')
// (17, 26, 'sp4_v_b_25')
// (17, 27, 'sp4_v_b_12')
// (17, 28, 'sp4_v_b_1')
// (18, 16, 'neigh_op_tnl_6')
// (18, 17, 'neigh_op_lft_6')
// (18, 18, 'neigh_op_bnl_6')

wire n1110;
// (16, 16, 'neigh_op_tnr_7')
// (16, 17, 'neigh_op_rgt_7')
// (16, 18, 'neigh_op_bnr_7')
// (17, 16, 'neigh_op_top_7')
// (17, 17, 'local_g2_7')
// (17, 17, 'lutff_6/in_3')
// (17, 17, 'lutff_7/out')
// (17, 18, 'neigh_op_bot_7')
// (18, 16, 'neigh_op_tnl_7')
// (18, 17, 'neigh_op_lft_7')
// (18, 18, 'neigh_op_bnl_7')

reg n1111 = 0;
// (16, 16, 'sp4_h_r_1')
// (17, 16, 'local_g1_4')
// (17, 16, 'lutff_2/in_3')
// (17, 16, 'sp4_h_r_12')
// (18, 16, 'sp4_h_r_25')
// (19, 16, 'sp4_h_r_36')
// (20, 16, 'sp4_h_l_36')
// (20, 16, 'sp4_h_r_1')
// (21, 16, 'sp4_h_r_12')
// (22, 16, 'sp4_h_r_25')
// (23, 12, 'neigh_op_tnr_2')
// (23, 13, 'neigh_op_rgt_2')
// (23, 13, 'sp4_r_v_b_36')
// (23, 14, 'neigh_op_bnr_2')
// (23, 14, 'sp4_r_v_b_25')
// (23, 15, 'sp4_r_v_b_12')
// (23, 16, 'sp4_h_r_36')
// (23, 16, 'sp4_r_v_b_1')
// (24, 12, 'neigh_op_top_2')
// (24, 12, 'sp4_v_t_36')
// (24, 13, 'lutff_2/out')
// (24, 13, 'sp4_v_b_36')
// (24, 14, 'neigh_op_bot_2')
// (24, 14, 'sp4_v_b_25')
// (24, 15, 'sp4_v_b_12')
// (24, 16, 'sp4_h_l_36')
// (24, 16, 'sp4_v_b_1')
// (25, 12, 'neigh_op_tnl_2')
// (25, 13, 'neigh_op_lft_2')
// (25, 14, 'neigh_op_bnl_2')

wire n1112;
// (16, 17, 'sp4_h_r_2')
// (17, 17, 'sp4_h_r_15')
// (18, 17, 'sp4_h_r_26')
// (19, 17, 'local_g2_7')
// (19, 17, 'lutff_4/in_3')
// (19, 17, 'sp4_h_r_39')
// (19, 18, 'sp4_r_v_b_45')
// (19, 19, 'sp4_r_v_b_32')
// (19, 20, 'neigh_op_tnr_4')
// (19, 20, 'sp4_r_v_b_21')
// (19, 21, 'neigh_op_rgt_4')
// (19, 21, 'sp4_r_v_b_8')
// (19, 22, 'neigh_op_bnr_4')
// (20, 17, 'sp4_h_l_39')
// (20, 17, 'sp4_v_t_45')
// (20, 18, 'sp4_v_b_45')
// (20, 19, 'sp4_v_b_32')
// (20, 20, 'neigh_op_top_4')
// (20, 20, 'sp4_v_b_21')
// (20, 21, 'lutff_4/out')
// (20, 21, 'sp4_v_b_8')
// (20, 22, 'neigh_op_bot_4')
// (21, 20, 'neigh_op_tnl_4')
// (21, 21, 'neigh_op_lft_4')
// (21, 22, 'neigh_op_bnl_4')

reg n1113 = 0;
// (16, 17, 'sp4_h_r_3')
// (17, 17, 'sp4_h_r_14')
// (18, 17, 'local_g3_3')
// (18, 17, 'lutff_7/in_1')
// (18, 17, 'sp4_h_r_27')
// (19, 17, 'sp4_h_r_38')
// (19, 18, 'sp4_r_v_b_38')
// (19, 19, 'sp4_r_v_b_27')
// (19, 20, 'sp4_r_v_b_14')
// (19, 21, 'sp4_r_v_b_3')
// (19, 22, 'sp4_r_v_b_37')
// (19, 23, 'sp4_r_v_b_24')
// (19, 24, 'neigh_op_tnr_0')
// (19, 24, 'sp4_r_v_b_13')
// (19, 25, 'neigh_op_rgt_0')
// (19, 25, 'sp4_r_v_b_0')
// (19, 26, 'neigh_op_bnr_0')
// (20, 17, 'sp4_h_l_38')
// (20, 17, 'sp4_v_t_38')
// (20, 18, 'sp4_v_b_38')
// (20, 19, 'sp4_v_b_27')
// (20, 20, 'sp4_v_b_14')
// (20, 21, 'sp4_v_b_3')
// (20, 21, 'sp4_v_t_37')
// (20, 22, 'sp4_v_b_37')
// (20, 23, 'sp4_v_b_24')
// (20, 24, 'neigh_op_top_0')
// (20, 24, 'sp4_v_b_13')
// (20, 25, 'lutff_0/out')
// (20, 25, 'sp4_v_b_0')
// (20, 26, 'neigh_op_bot_0')
// (21, 24, 'neigh_op_tnl_0')
// (21, 25, 'neigh_op_lft_0')
// (21, 26, 'neigh_op_bnl_0')

reg n1114 = 0;
// (16, 17, 'sp4_h_r_5')
// (17, 17, 'sp4_h_r_16')
// (18, 17, 'local_g2_5')
// (18, 17, 'lutff_4/in_1')
// (18, 17, 'sp4_h_r_29')
// (19, 17, 'sp4_h_r_40')
// (19, 18, 'sp4_r_v_b_40')
// (19, 19, 'neigh_op_tnr_0')
// (19, 19, 'sp4_r_v_b_29')
// (19, 20, 'neigh_op_rgt_0')
// (19, 20, 'sp4_r_v_b_16')
// (19, 21, 'neigh_op_bnr_0')
// (19, 21, 'sp4_r_v_b_5')
// (20, 17, 'sp4_h_l_40')
// (20, 17, 'sp4_v_t_40')
// (20, 18, 'sp4_v_b_40')
// (20, 19, 'neigh_op_top_0')
// (20, 19, 'sp4_v_b_29')
// (20, 20, 'lutff_0/out')
// (20, 20, 'sp4_v_b_16')
// (20, 21, 'neigh_op_bot_0')
// (20, 21, 'sp4_v_b_5')
// (21, 19, 'neigh_op_tnl_0')
// (21, 20, 'neigh_op_lft_0')
// (21, 21, 'neigh_op_bnl_0')

reg n1115 = 0;
// (16, 17, 'sp4_h_r_6')
// (17, 17, 'sp4_h_r_19')
// (18, 17, 'local_g3_6')
// (18, 17, 'lutff_0/in_3')
// (18, 17, 'sp4_h_r_30')
// (19, 17, 'sp4_h_r_43')
// (19, 18, 'neigh_op_tnr_7')
// (19, 18, 'sp4_r_v_b_43')
// (19, 19, 'neigh_op_rgt_7')
// (19, 19, 'sp4_r_v_b_30')
// (19, 20, 'neigh_op_bnr_7')
// (19, 20, 'sp4_r_v_b_19')
// (19, 21, 'sp4_r_v_b_6')
// (20, 17, 'sp4_h_l_43')
// (20, 17, 'sp4_v_t_43')
// (20, 18, 'neigh_op_top_7')
// (20, 18, 'sp4_v_b_43')
// (20, 19, 'lutff_7/out')
// (20, 19, 'sp4_v_b_30')
// (20, 20, 'neigh_op_bot_7')
// (20, 20, 'sp4_v_b_19')
// (20, 21, 'sp4_v_b_6')
// (21, 18, 'neigh_op_tnl_7')
// (21, 19, 'neigh_op_lft_7')
// (21, 20, 'neigh_op_bnl_7')

reg n1116 = 0;
// (16, 18, 'sp4_h_r_1')
// (17, 18, 'sp4_h_r_12')
// (18, 18, 'local_g2_1')
// (18, 18, 'lutff_0/in_3')
// (18, 18, 'sp4_h_r_25')
// (19, 18, 'neigh_op_tnr_5')
// (19, 18, 'sp4_h_r_36')
// (19, 19, 'neigh_op_rgt_5')
// (19, 19, 'sp4_r_v_b_42')
// (19, 20, 'neigh_op_bnr_5')
// (19, 20, 'sp4_r_v_b_31')
// (19, 21, 'sp4_r_v_b_18')
// (19, 22, 'sp4_r_v_b_7')
// (20, 18, 'neigh_op_top_5')
// (20, 18, 'sp4_h_l_36')
// (20, 18, 'sp4_v_t_42')
// (20, 19, 'lutff_5/out')
// (20, 19, 'sp4_v_b_42')
// (20, 20, 'neigh_op_bot_5')
// (20, 20, 'sp4_v_b_31')
// (20, 21, 'sp4_v_b_18')
// (20, 22, 'sp4_v_b_7')
// (21, 18, 'neigh_op_tnl_5')
// (21, 19, 'neigh_op_lft_5')
// (21, 20, 'neigh_op_bnl_5')

wire n1117;
// (16, 18, 'sp4_h_r_10')
// (17, 16, 'sp4_r_v_b_39')
// (17, 17, 'sp4_h_r_3')
// (17, 17, 'sp4_h_r_7')
// (17, 17, 'sp4_r_v_b_26')
// (17, 18, 'sp4_h_r_23')
// (17, 18, 'sp4_r_v_b_15')
// (17, 19, 'sp4_r_v_b_2')
// (18, 15, 'sp4_h_r_2')
// (18, 15, 'sp4_v_t_39')
// (18, 16, 'sp4_v_b_39')
// (18, 17, 'local_g0_2')
// (18, 17, 'lutff_global/cen')
// (18, 17, 'sp4_h_r_14')
// (18, 17, 'sp4_h_r_18')
// (18, 17, 'sp4_v_b_26')
// (18, 18, 'local_g2_2')
// (18, 18, 'lutff_global/cen')
// (18, 18, 'sp4_h_r_34')
// (18, 18, 'sp4_v_b_15')
// (18, 19, 'local_g0_2')
// (18, 19, 'lutff_global/cen')
// (18, 19, 'sp4_v_b_2')
// (19, 14, 'neigh_op_tnr_5')
// (19, 15, 'neigh_op_rgt_5')
// (19, 15, 'sp4_h_r_15')
// (19, 15, 'sp4_r_v_b_42')
// (19, 16, 'neigh_op_bnr_5')
// (19, 16, 'sp4_r_v_b_31')
// (19, 17, 'sp4_h_r_27')
// (19, 17, 'sp4_h_r_31')
// (19, 17, 'sp4_r_v_b_18')
// (19, 18, 'sp4_h_r_47')
// (19, 18, 'sp4_r_v_b_7')
// (20, 14, 'neigh_op_top_5')
// (20, 14, 'sp4_r_v_b_38')
// (20, 14, 'sp4_v_t_42')
// (20, 15, 'lutff_5/out')
// (20, 15, 'sp4_h_r_26')
// (20, 15, 'sp4_r_v_b_27')
// (20, 15, 'sp4_v_b_42')
// (20, 16, 'neigh_op_bot_5')
// (20, 16, 'sp4_r_v_b_14')
// (20, 16, 'sp4_v_b_31')
// (20, 17, 'sp4_h_r_38')
// (20, 17, 'sp4_h_r_42')
// (20, 17, 'sp4_r_v_b_3')
// (20, 17, 'sp4_v_b_18')
// (20, 18, 'sp4_h_l_47')
// (20, 18, 'sp4_h_r_7')
// (20, 18, 'sp4_v_b_7')
// (21, 13, 'sp4_v_t_38')
// (21, 14, 'neigh_op_tnl_5')
// (21, 14, 'sp4_v_b_38')
// (21, 15, 'neigh_op_lft_5')
// (21, 15, 'sp4_h_r_39')
// (21, 15, 'sp4_v_b_27')
// (21, 16, 'neigh_op_bnl_5')
// (21, 16, 'sp4_r_v_b_42')
// (21, 16, 'sp4_v_b_14')
// (21, 17, 'sp4_h_l_38')
// (21, 17, 'sp4_h_l_42')
// (21, 17, 'sp4_h_r_11')
// (21, 17, 'sp4_r_v_b_31')
// (21, 17, 'sp4_v_b_3')
// (21, 18, 'sp4_h_r_18')
// (21, 18, 'sp4_r_v_b_18')
// (21, 19, 'sp4_r_v_b_7')
// (21, 20, 'sp4_r_v_b_42')
// (21, 21, 'sp4_r_v_b_31')
// (21, 22, 'sp4_r_v_b_18')
// (21, 23, 'sp4_r_v_b_7')
// (22, 15, 'sp4_h_l_39')
// (22, 15, 'sp4_v_t_42')
// (22, 16, 'sp4_v_b_42')
// (22, 17, 'sp4_h_r_22')
// (22, 17, 'sp4_v_b_31')
// (22, 18, 'sp4_h_r_31')
// (22, 18, 'sp4_v_b_18')
// (22, 19, 'sp4_v_b_7')
// (22, 19, 'sp4_v_t_42')
// (22, 20, 'local_g2_2')
// (22, 20, 'lutff_global/cen')
// (22, 20, 'sp4_v_b_42')
// (22, 21, 'sp4_v_b_31')
// (22, 22, 'sp4_v_b_18')
// (22, 23, 'sp4_v_b_7')
// (23, 17, 'sp4_h_r_35')
// (23, 18, 'local_g2_2')
// (23, 18, 'lutff_global/cen')
// (23, 18, 'sp4_h_r_42')
// (24, 17, 'sp4_h_r_46')
// (24, 18, 'sp4_h_l_42')
// (25, 17, 'sp4_h_l_46')

reg n1118 = 0;
// (16, 18, 'sp4_h_r_4')
// (17, 18, 'sp4_h_r_17')
// (18, 18, 'local_g2_4')
// (18, 18, 'lutff_5/in_1')
// (18, 18, 'sp4_h_r_28')
// (19, 18, 'sp4_h_r_41')
// (19, 19, 'neigh_op_tnr_6')
// (19, 19, 'sp4_r_v_b_41')
// (19, 20, 'neigh_op_rgt_6')
// (19, 20, 'sp4_r_v_b_28')
// (19, 21, 'neigh_op_bnr_6')
// (19, 21, 'sp4_r_v_b_17')
// (19, 22, 'sp4_r_v_b_4')
// (20, 18, 'sp4_h_l_41')
// (20, 18, 'sp4_v_t_41')
// (20, 19, 'neigh_op_top_6')
// (20, 19, 'sp4_v_b_41')
// (20, 20, 'lutff_6/out')
// (20, 20, 'sp4_v_b_28')
// (20, 21, 'neigh_op_bot_6')
// (20, 21, 'sp4_v_b_17')
// (20, 22, 'sp4_v_b_4')
// (21, 19, 'neigh_op_tnl_6')
// (21, 20, 'neigh_op_lft_6')
// (21, 21, 'neigh_op_bnl_6')

wire n1119;
// (16, 19, 'neigh_op_tnr_0')
// (16, 20, 'neigh_op_rgt_0')
// (16, 21, 'neigh_op_bnr_0')
// (17, 19, 'neigh_op_top_0')
// (17, 20, 'local_g3_0')
// (17, 20, 'lutff_0/in_1')
// (17, 20, 'lutff_0/out')
// (17, 21, 'neigh_op_bot_0')
// (18, 19, 'neigh_op_tnl_0')
// (18, 20, 'neigh_op_lft_0')
// (18, 21, 'neigh_op_bnl_0')

wire n1120;
// (16, 19, 'neigh_op_tnr_1')
// (16, 20, 'neigh_op_rgt_1')
// (16, 21, 'neigh_op_bnr_1')
// (17, 19, 'neigh_op_top_1')
// (17, 20, 'local_g3_1')
// (17, 20, 'lutff_1/in_1')
// (17, 20, 'lutff_1/out')
// (17, 21, 'neigh_op_bot_1')
// (18, 19, 'neigh_op_tnl_1')
// (18, 20, 'neigh_op_lft_1')
// (18, 21, 'neigh_op_bnl_1')

wire n1121;
// (16, 19, 'neigh_op_tnr_2')
// (16, 20, 'neigh_op_rgt_2')
// (16, 21, 'neigh_op_bnr_2')
// (17, 19, 'neigh_op_top_2')
// (17, 20, 'local_g1_2')
// (17, 20, 'lutff_2/in_1')
// (17, 20, 'lutff_2/out')
// (17, 21, 'neigh_op_bot_2')
// (18, 19, 'neigh_op_tnl_2')
// (18, 20, 'neigh_op_lft_2')
// (18, 21, 'neigh_op_bnl_2')

wire n1122;
// (16, 19, 'neigh_op_tnr_3')
// (16, 20, 'neigh_op_rgt_3')
// (16, 21, 'neigh_op_bnr_3')
// (17, 19, 'neigh_op_top_3')
// (17, 20, 'local_g1_3')
// (17, 20, 'lutff_3/in_1')
// (17, 20, 'lutff_3/out')
// (17, 21, 'neigh_op_bot_3')
// (18, 19, 'neigh_op_tnl_3')
// (18, 20, 'neigh_op_lft_3')
// (18, 21, 'neigh_op_bnl_3')

wire n1123;
// (16, 19, 'neigh_op_tnr_4')
// (16, 20, 'neigh_op_rgt_4')
// (16, 21, 'neigh_op_bnr_4')
// (17, 19, 'neigh_op_top_4')
// (17, 20, 'local_g3_4')
// (17, 20, 'lutff_4/in_1')
// (17, 20, 'lutff_4/out')
// (17, 21, 'neigh_op_bot_4')
// (18, 19, 'neigh_op_tnl_4')
// (18, 20, 'neigh_op_lft_4')
// (18, 21, 'neigh_op_bnl_4')

wire n1124;
// (16, 19, 'neigh_op_tnr_5')
// (16, 20, 'neigh_op_rgt_5')
// (16, 21, 'neigh_op_bnr_5')
// (17, 19, 'neigh_op_top_5')
// (17, 20, 'local_g1_5')
// (17, 20, 'lutff_5/in_1')
// (17, 20, 'lutff_5/out')
// (17, 21, 'neigh_op_bot_5')
// (18, 19, 'neigh_op_tnl_5')
// (18, 20, 'neigh_op_lft_5')
// (18, 21, 'neigh_op_bnl_5')

wire n1125;
// (16, 19, 'neigh_op_tnr_6')
// (16, 20, 'neigh_op_rgt_6')
// (16, 21, 'neigh_op_bnr_6')
// (17, 19, 'neigh_op_top_6')
// (17, 20, 'local_g1_6')
// (17, 20, 'lutff_6/in_1')
// (17, 20, 'lutff_6/out')
// (17, 21, 'neigh_op_bot_6')
// (18, 19, 'neigh_op_tnl_6')
// (18, 20, 'neigh_op_lft_6')
// (18, 21, 'neigh_op_bnl_6')

wire n1126;
// (16, 19, 'neigh_op_tnr_7')
// (16, 20, 'neigh_op_rgt_7')
// (16, 21, 'neigh_op_bnr_7')
// (17, 19, 'neigh_op_top_7')
// (17, 20, 'local_g1_7')
// (17, 20, 'lutff_7/in_1')
// (17, 20, 'lutff_7/out')
// (17, 21, 'neigh_op_bot_7')
// (18, 19, 'neigh_op_tnl_7')
// (18, 20, 'neigh_op_lft_7')
// (18, 21, 'neigh_op_bnl_7')

wire n1127;
// (16, 19, 'sp4_r_v_b_40')
// (16, 20, 'neigh_op_tnr_0')
// (16, 20, 'sp4_r_v_b_29')
// (16, 21, 'neigh_op_rgt_0')
// (16, 21, 'sp4_r_v_b_16')
// (16, 22, 'local_g0_0')
// (16, 22, 'local_g1_0')
// (16, 22, 'lutff_0/in_3')
// (16, 22, 'lutff_1/in_1')
// (16, 22, 'lutff_2/in_3')
// (16, 22, 'lutff_3/in_1')
// (16, 22, 'lutff_4/in_2')
// (16, 22, 'neigh_op_bnr_0')
// (16, 22, 'sp4_r_v_b_5')
// (17, 18, 'sp4_v_t_40')
// (17, 19, 'sp4_v_b_40')
// (17, 20, 'neigh_op_top_0')
// (17, 20, 'sp4_r_v_b_44')
// (17, 20, 'sp4_v_b_29')
// (17, 21, 'lutff_0/out')
// (17, 21, 'sp4_r_v_b_33')
// (17, 21, 'sp4_v_b_16')
// (17, 22, 'neigh_op_bot_0')
// (17, 22, 'sp4_h_r_5')
// (17, 22, 'sp4_r_v_b_20')
// (17, 22, 'sp4_v_b_5')
// (17, 23, 'sp4_r_v_b_9')
// (18, 19, 'sp4_v_t_44')
// (18, 20, 'neigh_op_tnl_0')
// (18, 20, 'sp4_v_b_44')
// (18, 21, 'local_g0_0')
// (18, 21, 'local_g1_0')
// (18, 21, 'lutff_0/in_2')
// (18, 21, 'lutff_1/in_2')
// (18, 21, 'lutff_2/in_0')
// (18, 21, 'lutff_3/in_2')
// (18, 21, 'lutff_4/in_1')
// (18, 21, 'lutff_5/in_2')
// (18, 21, 'lutff_6/in_1')
// (18, 21, 'lutff_7/in_2')
// (18, 21, 'neigh_op_lft_0')
// (18, 21, 'sp4_v_b_33')
// (18, 22, 'local_g2_0')
// (18, 22, 'lutff_2/in_2')
// (18, 22, 'neigh_op_bnl_0')
// (18, 22, 'sp4_h_r_16')
// (18, 22, 'sp4_v_b_20')
// (18, 23, 'local_g0_1')
// (18, 23, 'local_g1_1')
// (18, 23, 'lutff_0/in_1')
// (18, 23, 'lutff_1/in_2')
// (18, 23, 'lutff_2/in_2')
// (18, 23, 'lutff_3/in_2')
// (18, 23, 'lutff_4/in_1')
// (18, 23, 'lutff_5/in_2')
// (18, 23, 'lutff_6/in_1')
// (18, 23, 'lutff_7/in_2')
// (18, 23, 'sp4_v_b_9')
// (19, 22, 'sp4_h_r_29')
// (20, 22, 'local_g2_0')
// (20, 22, 'local_g3_0')
// (20, 22, 'lutff_5/in_3')
// (20, 22, 'lutff_6/in_1')
// (20, 22, 'sp4_h_r_40')
// (21, 22, 'sp4_h_l_40')

wire n1128;
// (16, 20, 'neigh_op_tnr_5')
// (16, 21, 'neigh_op_rgt_5')
// (16, 22, 'neigh_op_bnr_5')
// (17, 20, 'neigh_op_top_5')
// (17, 21, 'lutff_5/out')
// (17, 22, 'neigh_op_bot_5')
// (18, 20, 'local_g3_5')
// (18, 20, 'lutff_7/in_3')
// (18, 20, 'neigh_op_tnl_5')
// (18, 21, 'neigh_op_lft_5')
// (18, 22, 'neigh_op_bnl_5')

wire n1129;
// (16, 21, 'neigh_op_tnr_0')
// (16, 22, 'neigh_op_rgt_0')
// (16, 23, 'neigh_op_bnr_0')
// (17, 21, 'neigh_op_top_0')
// (17, 22, 'local_g3_0')
// (17, 22, 'lutff_0/in_1')
// (17, 22, 'lutff_0/out')
// (17, 23, 'neigh_op_bot_0')
// (18, 21, 'neigh_op_tnl_0')
// (18, 22, 'neigh_op_lft_0')
// (18, 23, 'neigh_op_bnl_0')

wire n1130;
// (16, 21, 'neigh_op_tnr_1')
// (16, 22, 'neigh_op_rgt_1')
// (16, 23, 'neigh_op_bnr_1')
// (17, 21, 'neigh_op_top_1')
// (17, 22, 'local_g1_1')
// (17, 22, 'lutff_1/in_1')
// (17, 22, 'lutff_1/out')
// (17, 23, 'neigh_op_bot_1')
// (18, 21, 'neigh_op_tnl_1')
// (18, 22, 'neigh_op_lft_1')
// (18, 23, 'neigh_op_bnl_1')

wire n1131;
// (16, 21, 'neigh_op_tnr_2')
// (16, 22, 'neigh_op_rgt_2')
// (16, 23, 'neigh_op_bnr_2')
// (17, 21, 'neigh_op_top_2')
// (17, 22, 'local_g0_2')
// (17, 22, 'lutff_2/in_2')
// (17, 22, 'lutff_2/out')
// (17, 23, 'neigh_op_bot_2')
// (18, 21, 'neigh_op_tnl_2')
// (18, 22, 'neigh_op_lft_2')
// (18, 23, 'neigh_op_bnl_2')

wire n1132;
// (16, 21, 'neigh_op_tnr_3')
// (16, 22, 'neigh_op_rgt_3')
// (16, 23, 'neigh_op_bnr_3')
// (17, 21, 'neigh_op_top_3')
// (17, 22, 'local_g2_3')
// (17, 22, 'lutff_3/in_2')
// (17, 22, 'lutff_3/out')
// (17, 23, 'neigh_op_bot_3')
// (18, 21, 'neigh_op_tnl_3')
// (18, 22, 'neigh_op_lft_3')
// (18, 23, 'neigh_op_bnl_3')

wire n1133;
// (16, 21, 'neigh_op_tnr_4')
// (16, 22, 'neigh_op_rgt_4')
// (16, 23, 'neigh_op_bnr_4')
// (17, 21, 'neigh_op_top_4')
// (17, 22, 'local_g0_4')
// (17, 22, 'lutff_4/in_2')
// (17, 22, 'lutff_4/out')
// (17, 23, 'neigh_op_bot_4')
// (18, 21, 'neigh_op_tnl_4')
// (18, 22, 'neigh_op_lft_4')
// (18, 23, 'neigh_op_bnl_4')

wire n1134;
// (16, 21, 'neigh_op_tnr_5')
// (16, 22, 'neigh_op_rgt_5')
// (16, 23, 'neigh_op_bnr_5')
// (17, 21, 'neigh_op_top_5')
// (17, 22, 'local_g0_5')
// (17, 22, 'lutff_5/in_2')
// (17, 22, 'lutff_5/out')
// (17, 23, 'neigh_op_bot_5')
// (18, 21, 'neigh_op_tnl_5')
// (18, 22, 'neigh_op_lft_5')
// (18, 23, 'neigh_op_bnl_5')

wire n1135;
// (16, 21, 'neigh_op_tnr_6')
// (16, 22, 'neigh_op_rgt_6')
// (16, 23, 'neigh_op_bnr_6')
// (17, 21, 'neigh_op_top_6')
// (17, 22, 'local_g2_6')
// (17, 22, 'lutff_6/in_2')
// (17, 22, 'lutff_6/out')
// (17, 23, 'neigh_op_bot_6')
// (18, 21, 'neigh_op_tnl_6')
// (18, 22, 'neigh_op_lft_6')
// (18, 23, 'neigh_op_bnl_6')

wire n1136;
// (16, 21, 'neigh_op_tnr_7')
// (16, 22, 'neigh_op_rgt_7')
// (16, 23, 'neigh_op_bnr_7')
// (17, 21, 'neigh_op_top_7')
// (17, 22, 'local_g0_7')
// (17, 22, 'lutff_7/in_2')
// (17, 22, 'lutff_7/out')
// (17, 23, 'neigh_op_bot_7')
// (18, 21, 'neigh_op_tnl_7')
// (18, 22, 'neigh_op_lft_7')
// (18, 23, 'neigh_op_bnl_7')

wire n1137;
// (16, 22, 'neigh_op_tnr_0')
// (16, 23, 'neigh_op_rgt_0')
// (16, 24, 'neigh_op_bnr_0')
// (17, 22, 'neigh_op_top_0')
// (17, 23, 'local_g2_0')
// (17, 23, 'lutff_0/in_2')
// (17, 23, 'lutff_0/out')
// (17, 24, 'neigh_op_bot_0')
// (18, 22, 'neigh_op_tnl_0')
// (18, 23, 'neigh_op_lft_0')
// (18, 24, 'neigh_op_bnl_0')

wire n1138;
// (16, 22, 'neigh_op_tnr_1')
// (16, 23, 'neigh_op_rgt_1')
// (16, 24, 'neigh_op_bnr_1')
// (17, 22, 'neigh_op_top_1')
// (17, 23, 'local_g1_2')
// (17, 23, 'lutff_1/in_2')
// (17, 23, 'lutff_1/out')
// (17, 23, 'sp4_h_r_2')
// (17, 24, 'neigh_op_bot_1')
// (18, 22, 'neigh_op_tnl_1')
// (18, 23, 'neigh_op_lft_1')
// (18, 23, 'sp4_h_r_15')
// (18, 24, 'neigh_op_bnl_1')
// (19, 23, 'sp4_h_r_26')
// (20, 23, 'sp4_h_r_39')
// (21, 23, 'sp4_h_l_39')

wire n1139;
// (16, 22, 'neigh_op_tnr_2')
// (16, 23, 'neigh_op_rgt_2')
// (16, 24, 'neigh_op_bnr_2')
// (17, 22, 'neigh_op_top_2')
// (17, 23, 'local_g0_2')
// (17, 23, 'lutff_2/in_2')
// (17, 23, 'lutff_2/out')
// (17, 24, 'neigh_op_bot_2')
// (18, 22, 'neigh_op_tnl_2')
// (18, 23, 'neigh_op_lft_2')
// (18, 24, 'neigh_op_bnl_2')

wire n1140;
// (16, 22, 'neigh_op_tnr_3')
// (16, 23, 'neigh_op_rgt_3')
// (16, 24, 'neigh_op_bnr_3')
// (17, 22, 'neigh_op_top_3')
// (17, 23, 'local_g3_3')
// (17, 23, 'lutff_3/in_1')
// (17, 23, 'lutff_3/out')
// (17, 24, 'neigh_op_bot_3')
// (18, 22, 'neigh_op_tnl_3')
// (18, 23, 'neigh_op_lft_3')
// (18, 24, 'neigh_op_bnl_3')

wire n1141;
// (16, 22, 'neigh_op_tnr_4')
// (16, 23, 'neigh_op_rgt_4')
// (16, 24, 'neigh_op_bnr_4')
// (17, 22, 'neigh_op_top_4')
// (17, 23, 'local_g0_4')
// (17, 23, 'lutff_4/in_2')
// (17, 23, 'lutff_4/out')
// (17, 24, 'neigh_op_bot_4')
// (18, 22, 'neigh_op_tnl_4')
// (18, 23, 'neigh_op_lft_4')
// (18, 24, 'neigh_op_bnl_4')

wire n1142;
// (16, 22, 'neigh_op_tnr_5')
// (16, 23, 'neigh_op_rgt_5')
// (16, 24, 'neigh_op_bnr_5')
// (17, 22, 'neigh_op_top_5')
// (17, 23, 'local_g0_5')
// (17, 23, 'lutff_5/in_2')
// (17, 23, 'lutff_5/out')
// (17, 24, 'neigh_op_bot_5')
// (18, 22, 'neigh_op_tnl_5')
// (18, 23, 'neigh_op_lft_5')
// (18, 24, 'neigh_op_bnl_5')

wire n1143;
// (16, 22, 'neigh_op_tnr_6')
// (16, 23, 'neigh_op_rgt_6')
// (16, 24, 'neigh_op_bnr_6')
// (17, 22, 'neigh_op_top_6')
// (17, 23, 'local_g2_6')
// (17, 23, 'lutff_6/in_2')
// (17, 23, 'lutff_6/out')
// (17, 24, 'neigh_op_bot_6')
// (18, 22, 'neigh_op_tnl_6')
// (18, 23, 'neigh_op_lft_6')
// (18, 24, 'neigh_op_bnl_6')

wire n1144;
// (16, 22, 'neigh_op_tnr_7')
// (16, 23, 'neigh_op_rgt_7')
// (16, 24, 'neigh_op_bnr_7')
// (17, 22, 'neigh_op_top_7')
// (17, 23, 'local_g2_7')
// (17, 23, 'lutff_7/in_2')
// (17, 23, 'lutff_7/out')
// (17, 24, 'neigh_op_bot_7')
// (18, 22, 'neigh_op_tnl_7')
// (18, 23, 'neigh_op_lft_7')
// (18, 24, 'neigh_op_bnl_7')

wire n1145;
// (16, 22, 'sp4_h_r_0')
// (17, 21, 'neigh_op_tnr_4')
// (17, 22, 'neigh_op_rgt_4')
// (17, 22, 'sp4_h_r_13')
// (17, 23, 'neigh_op_bnr_4')
// (18, 21, 'neigh_op_top_4')
// (18, 22, 'lutff_4/out')
// (18, 22, 'sp4_h_r_24')
// (18, 23, 'neigh_op_bot_4')
// (19, 19, 'sp4_r_v_b_43')
// (19, 20, 'sp4_r_v_b_30')
// (19, 21, 'local_g3_3')
// (19, 21, 'lutff_global/cen')
// (19, 21, 'neigh_op_tnl_4')
// (19, 21, 'sp4_r_v_b_19')
// (19, 22, 'neigh_op_lft_4')
// (19, 22, 'sp4_h_r_37')
// (19, 22, 'sp4_r_v_b_6')
// (19, 23, 'neigh_op_bnl_4')
// (20, 18, 'sp4_v_t_43')
// (20, 19, 'sp4_v_b_43')
// (20, 20, 'sp4_v_b_30')
// (20, 21, 'sp4_v_b_19')
// (20, 22, 'sp4_h_l_37')
// (20, 22, 'sp4_v_b_6')

wire n1146;
// (16, 22, 'sp4_r_v_b_43')
// (16, 23, 'sp4_r_v_b_30')
// (16, 24, 'sp4_r_v_b_19')
// (16, 25, 'sp4_r_v_b_6')
// (17, 19, 'sp12_v_t_23')
// (17, 20, 'sp12_v_b_23')
// (17, 21, 'sp12_v_b_20')
// (17, 21, 'sp4_h_r_6')
// (17, 21, 'sp4_v_t_43')
// (17, 22, 'sp12_v_b_19')
// (17, 22, 'sp4_v_b_43')
// (17, 23, 'sp12_v_b_16')
// (17, 23, 'sp4_v_b_30')
// (17, 24, 'sp12_v_b_15')
// (17, 24, 'sp4_v_b_19')
// (17, 25, 'sp12_v_b_12')
// (17, 25, 'sp4_v_b_6')
// (17, 26, 'sp12_v_b_11')
// (17, 27, 'sp12_v_b_8')
// (17, 28, 'sp12_v_b_7')
// (17, 29, 'sp12_v_b_4')
// (17, 30, 'sp12_v_b_3')
// (17, 31, 'sp12_h_r_0')
// (17, 31, 'sp12_v_b_0')
// (18, 21, 'sp4_h_r_19')
// (18, 31, 'sp12_h_r_3')
// (19, 21, 'local_g2_6')
// (19, 21, 'lutff_3/in_1')
// (19, 21, 'sp4_h_r_30')
// (19, 31, 'sp12_h_r_4')
// (20, 21, 'sp4_h_r_43')
// (20, 31, 'sp12_h_r_7')
// (21, 21, 'sp4_h_l_43')
// (21, 31, 'sp12_h_r_8')
// (22, 31, 'sp12_h_r_11')
// (23, 31, 'sp12_h_r_12')
// (24, 31, 'sp12_h_r_15')
// (25, 31, 'sp12_h_r_16')
// (26, 31, 'sp12_h_r_19')
// (27, 31, 'sp12_h_r_20')
// (28, 31, 'sp12_h_r_23')
// (28, 32, 'neigh_op_tnr_2')
// (28, 32, 'neigh_op_tnr_6')
// (29, 31, 'sp12_h_l_23')
// (29, 31, 'sp12_v_t_23')
// (29, 32, 'neigh_op_top_2')
// (29, 32, 'neigh_op_top_6')
// (29, 32, 'sp12_v_b_23')
// (29, 33, 'io_1/D_IN_0')
// (29, 33, 'span12_vert_20')
// (30, 32, 'neigh_op_tnl_2')
// (30, 32, 'neigh_op_tnl_6')

reg io_33_4_0 = 0;
// (16, 23, 'sp12_h_r_0')
// (17, 22, 'neigh_op_tnr_6')
// (17, 23, 'neigh_op_rgt_6')
// (17, 23, 'sp12_h_r_3')
// (17, 24, 'neigh_op_bnr_6')
// (18, 22, 'neigh_op_top_6')
// (18, 23, 'lutff_6/out')
// (18, 23, 'sp12_h_r_4')
// (18, 24, 'neigh_op_bot_6')
// (19, 22, 'neigh_op_tnl_6')
// (19, 23, 'neigh_op_lft_6')
// (19, 23, 'sp12_h_r_7')
// (19, 24, 'neigh_op_bnl_6')
// (20, 23, 'sp12_h_r_8')
// (21, 23, 'sp12_h_r_11')
// (22, 23, 'sp12_h_r_12')
// (23, 23, 'sp12_h_r_15')
// (24, 23, 'sp12_h_r_16')
// (25, 23, 'sp12_h_r_19')
// (26, 23, 'sp12_h_r_20')
// (27, 12, 'sp4_r_v_b_45')
// (27, 13, 'sp4_r_v_b_32')
// (27, 14, 'sp4_r_v_b_21')
// (27, 15, 'sp4_r_v_b_8')
// (27, 23, 'sp12_h_r_23')
// (28, 11, 'sp12_v_t_23')
// (28, 11, 'sp4_h_r_8')
// (28, 11, 'sp4_v_t_45')
// (28, 12, 'sp12_v_b_23')
// (28, 12, 'sp4_v_b_45')
// (28, 13, 'sp12_v_b_20')
// (28, 13, 'sp4_v_b_32')
// (28, 14, 'sp12_v_b_19')
// (28, 14, 'sp4_v_b_21')
// (28, 15, 'sp12_v_b_16')
// (28, 15, 'sp4_v_b_8')
// (28, 16, 'sp12_v_b_15')
// (28, 17, 'sp12_v_b_12')
// (28, 18, 'sp12_v_b_11')
// (28, 19, 'sp12_v_b_8')
// (28, 20, 'sp12_v_b_7')
// (28, 21, 'sp12_v_b_4')
// (28, 22, 'sp12_v_b_3')
// (28, 23, 'sp12_h_l_23')
// (28, 23, 'sp12_v_b_0')
// (29, 11, 'sp4_h_r_21')
// (30, 11, 'sp4_h_r_32')
// (31, 8, 'sp4_r_v_b_39')
// (31, 9, 'sp4_r_v_b_26')
// (31, 10, 'sp4_r_v_b_15')
// (31, 11, 'sp4_h_r_45')
// (31, 11, 'sp4_r_v_b_2')
// (32, 7, 'sp4_h_r_7')
// (32, 7, 'sp4_v_t_39')
// (32, 8, 'sp4_v_b_39')
// (32, 9, 'sp4_v_b_26')
// (32, 10, 'sp4_v_b_15')
// (32, 11, 'sp4_h_l_45')
// (32, 11, 'sp4_v_b_2')
// (33, 3, 'span4_vert_t_13')
// (33, 4, 'io_0/D_OUT_0')
// (33, 4, 'io_0/PAD')
// (33, 4, 'local_g1_5')
// (33, 4, 'span4_vert_b_13')
// (33, 5, 'span4_vert_b_9')
// (33, 6, 'span4_vert_b_5')
// (33, 7, 'span4_horz_7')
// (33, 7, 'span4_vert_b_1')

reg n1148 = 0;
// (16, 23, 'sp12_h_r_1')
// (17, 23, 'sp12_h_r_2')
// (18, 22, 'neigh_op_tnr_7')
// (18, 23, 'neigh_op_rgt_7')
// (18, 23, 'sp12_h_r_5')
// (18, 24, 'neigh_op_bnr_7')
// (19, 22, 'neigh_op_top_7')
// (19, 23, 'local_g2_7')
// (19, 23, 'lutff_7/in_2')
// (19, 23, 'lutff_7/out')
// (19, 23, 'sp12_h_r_6')
// (19, 24, 'neigh_op_bot_7')
// (20, 22, 'neigh_op_tnl_7')
// (20, 23, 'neigh_op_lft_7')
// (20, 23, 'sp12_h_r_9')
// (20, 24, 'neigh_op_bnl_7')
// (21, 23, 'sp12_h_r_10')
// (22, 23, 'sp12_h_r_13')
// (23, 23, 'sp12_h_r_14')
// (24, 23, 'sp12_h_r_17')
// (25, 23, 'sp12_h_r_18')
// (26, 23, 'sp12_h_r_21')
// (26, 23, 'sp4_h_r_10')
// (27, 23, 'sp12_h_r_22')
// (27, 23, 'sp4_h_r_23')
// (28, 23, 'sp12_h_l_22')
// (28, 23, 'sp4_h_r_34')
// (29, 16, 'sp4_r_v_b_37')
// (29, 17, 'sp4_r_v_b_24')
// (29, 18, 'sp4_r_v_b_13')
// (29, 19, 'sp4_r_v_b_0')
// (29, 20, 'sp4_r_v_b_41')
// (29, 21, 'sp4_r_v_b_28')
// (29, 22, 'sp4_r_v_b_17')
// (29, 23, 'sp4_h_r_47')
// (29, 23, 'sp4_r_v_b_4')
// (30, 15, 'sp4_h_r_5')
// (30, 15, 'sp4_v_t_37')
// (30, 16, 'sp4_v_b_37')
// (30, 17, 'sp4_v_b_24')
// (30, 18, 'sp4_v_b_13')
// (30, 19, 'sp4_v_b_0')
// (30, 19, 'sp4_v_t_41')
// (30, 20, 'sp4_v_b_41')
// (30, 21, 'sp4_v_b_28')
// (30, 22, 'sp4_v_b_17')
// (30, 23, 'sp4_h_l_47')
// (30, 23, 'sp4_v_b_4')
// (31, 15, 'sp4_h_r_16')
// (32, 15, 'sp4_h_r_29')
// (33, 15, 'io_1/OUT_ENB')
// (33, 15, 'local_g1_5')
// (33, 15, 'span4_horz_29')

wire n1149;
// (16, 24, 'neigh_op_tnr_3')
// (16, 25, 'neigh_op_rgt_3')
// (16, 26, 'neigh_op_bnr_3')
// (17, 22, 'sp4_r_v_b_42')
// (17, 23, 'sp4_r_v_b_31')
// (17, 24, 'neigh_op_top_3')
// (17, 24, 'sp4_r_v_b_18')
// (17, 25, 'lutff_3/out')
// (17, 25, 'sp4_r_v_b_7')
// (17, 26, 'neigh_op_bot_3')
// (18, 21, 'sp4_h_r_0')
// (18, 21, 'sp4_v_t_42')
// (18, 22, 'sp4_v_b_42')
// (18, 23, 'sp4_v_b_31')
// (18, 24, 'neigh_op_tnl_3')
// (18, 24, 'sp4_v_b_18')
// (18, 25, 'neigh_op_lft_3')
// (18, 25, 'sp4_v_b_7')
// (18, 26, 'neigh_op_bnl_3')
// (19, 21, 'sp4_h_r_13')
// (20, 21, 'sp4_h_r_24')
// (21, 21, 'local_g3_5')
// (21, 21, 'lutff_7/in_3')
// (21, 21, 'sp4_h_r_37')
// (22, 21, 'sp4_h_l_37')

reg n1150 = 0;
// (16, 24, 'sp4_r_v_b_37')
// (16, 25, 'sp4_r_v_b_24')
// (16, 26, 'sp4_r_v_b_13')
// (16, 27, 'sp4_r_v_b_0')
// (17, 23, 'sp4_h_r_0')
// (17, 23, 'sp4_v_t_37')
// (17, 24, 'sp4_v_b_37')
// (17, 25, 'local_g2_0')
// (17, 25, 'lutff_3/in_1')
// (17, 25, 'sp4_v_b_24')
// (17, 26, 'sp4_v_b_13')
// (17, 27, 'sp4_v_b_0')
// (18, 23, 'sp4_h_r_13')
// (19, 19, 'neigh_op_tnr_2')
// (19, 20, 'neigh_op_rgt_2')
// (19, 21, 'neigh_op_bnr_2')
// (19, 23, 'sp4_h_r_24')
// (20, 19, 'neigh_op_top_2')
// (20, 20, 'lutff_2/out')
// (20, 20, 'sp4_r_v_b_37')
// (20, 21, 'neigh_op_bot_2')
// (20, 21, 'sp4_r_v_b_24')
// (20, 22, 'sp4_r_v_b_13')
// (20, 23, 'sp4_h_r_37')
// (20, 23, 'sp4_r_v_b_0')
// (21, 19, 'neigh_op_tnl_2')
// (21, 19, 'sp4_v_t_37')
// (21, 20, 'neigh_op_lft_2')
// (21, 20, 'sp4_v_b_37')
// (21, 21, 'neigh_op_bnl_2')
// (21, 21, 'sp4_v_b_24')
// (21, 22, 'sp4_v_b_13')
// (21, 23, 'sp4_h_l_37')
// (21, 23, 'sp4_v_b_0')

reg n1151 = 0;
// (16, 25, 'sp4_h_r_1')
// (17, 25, 'sp4_h_r_12')
// (18, 25, 'local_g2_1')
// (18, 25, 'lutff_2/in_1')
// (18, 25, 'sp4_h_r_25')
// (19, 25, 'neigh_op_tnr_2')
// (19, 25, 'sp4_h_r_36')
// (19, 26, 'neigh_op_rgt_2')
// (19, 26, 'sp4_r_v_b_36')
// (19, 27, 'neigh_op_bnr_2')
// (19, 27, 'sp4_r_v_b_25')
// (19, 28, 'sp4_r_v_b_12')
// (19, 29, 'sp4_r_v_b_1')
// (20, 25, 'neigh_op_top_2')
// (20, 25, 'sp4_h_l_36')
// (20, 25, 'sp4_v_t_36')
// (20, 26, 'lutff_2/out')
// (20, 26, 'sp4_v_b_36')
// (20, 27, 'neigh_op_bot_2')
// (20, 27, 'sp4_v_b_25')
// (20, 28, 'sp4_v_b_12')
// (20, 29, 'sp4_v_b_1')
// (21, 25, 'neigh_op_tnl_2')
// (21, 26, 'neigh_op_lft_2')
// (21, 27, 'neigh_op_bnl_2')

reg n1152 = 0;
// (17, 4, 'sp12_v_t_23')
// (17, 5, 'sp12_v_b_23')
// (17, 6, 'sp12_v_b_20')
// (17, 7, 'sp12_v_b_19')
// (17, 8, 'sp12_v_b_16')
// (17, 9, 'sp12_v_b_15')
// (17, 10, 'sp12_v_b_12')
// (17, 11, 'sp12_v_b_11')
// (17, 12, 'local_g2_0')
// (17, 12, 'lutff_7/in_1')
// (17, 12, 'sp12_v_b_8')
// (17, 13, 'sp12_v_b_7')
// (17, 14, 'sp12_v_b_4')
// (17, 15, 'sp12_v_b_3')
// (17, 16, 'sp12_h_r_0')
// (17, 16, 'sp12_v_b_0')
// (18, 16, 'sp12_h_r_3')
// (19, 16, 'sp12_h_r_4')
// (20, 16, 'sp12_h_r_7')
// (21, 16, 'sp12_h_r_8')
// (22, 15, 'neigh_op_tnr_2')
// (22, 16, 'neigh_op_rgt_2')
// (22, 16, 'sp12_h_r_11')
// (22, 17, 'neigh_op_bnr_2')
// (23, 15, 'neigh_op_top_2')
// (23, 16, 'lutff_2/out')
// (23, 16, 'sp12_h_r_12')
// (23, 17, 'neigh_op_bot_2')
// (24, 15, 'neigh_op_tnl_2')
// (24, 16, 'neigh_op_lft_2')
// (24, 16, 'sp12_h_r_15')
// (24, 17, 'neigh_op_bnl_2')
// (25, 16, 'sp12_h_r_16')
// (26, 16, 'sp12_h_r_19')
// (27, 16, 'sp12_h_r_20')
// (28, 16, 'sp12_h_r_23')
// (29, 16, 'sp12_h_l_23')

reg n1153 = 0;
// (17, 7, 'sp12_v_t_23')
// (17, 8, 'sp12_v_b_23')
// (17, 9, 'sp12_v_b_20')
// (17, 10, 'sp12_v_b_19')
// (17, 11, 'sp12_v_b_16')
// (17, 12, 'sp12_v_b_15')
// (17, 13, 'sp12_v_b_12')
// (17, 14, 'sp12_v_b_11')
// (17, 15, 'local_g2_0')
// (17, 15, 'lutff_4/in_0')
// (17, 15, 'sp12_v_b_8')
// (17, 16, 'sp12_v_b_7')
// (17, 17, 'sp12_v_b_4')
// (17, 18, 'sp12_v_b_3')
// (17, 19, 'sp12_h_r_0')
// (17, 19, 'sp12_v_b_0')
// (18, 18, 'neigh_op_tnr_6')
// (18, 19, 'neigh_op_rgt_6')
// (18, 19, 'sp12_h_r_3')
// (18, 20, 'neigh_op_bnr_6')
// (19, 18, 'neigh_op_top_6')
// (19, 19, 'lutff_6/out')
// (19, 19, 'sp12_h_r_4')
// (19, 20, 'neigh_op_bot_6')
// (20, 18, 'neigh_op_tnl_6')
// (20, 19, 'neigh_op_lft_6')
// (20, 19, 'sp12_h_r_7')
// (20, 20, 'neigh_op_bnl_6')
// (21, 19, 'sp12_h_r_8')
// (22, 19, 'sp12_h_r_11')
// (23, 19, 'sp12_h_r_12')
// (24, 19, 'sp12_h_r_15')
// (25, 19, 'sp12_h_r_16')
// (26, 19, 'sp12_h_r_19')
// (27, 19, 'sp12_h_r_20')
// (28, 19, 'sp12_h_r_23')
// (29, 19, 'sp12_h_l_23')

reg n1154 = 0;
// (17, 7, 'sp4_r_v_b_46')
// (17, 8, 'neigh_op_tnr_3')
// (17, 8, 'sp4_r_v_b_35')
// (17, 9, 'neigh_op_rgt_3')
// (17, 9, 'sp4_r_v_b_22')
// (17, 10, 'neigh_op_bnr_3')
// (17, 10, 'sp4_r_v_b_11')
// (18, 6, 'sp4_v_t_46')
// (18, 7, 'local_g3_6')
// (18, 7, 'lutff_0/in_3')
// (18, 7, 'sp4_v_b_46')
// (18, 8, 'neigh_op_top_3')
// (18, 8, 'sp4_v_b_35')
// (18, 9, 'lutff_3/out')
// (18, 9, 'sp4_v_b_22')
// (18, 10, 'neigh_op_bot_3')
// (18, 10, 'sp4_v_b_11')
// (19, 8, 'neigh_op_tnl_3')
// (19, 9, 'neigh_op_lft_3')
// (19, 10, 'neigh_op_bnl_3')

reg n1155 = 0;
// (17, 8, 'local_g2_0')
// (17, 8, 'lutff_5/in_3')
// (17, 8, 'neigh_op_tnr_0')
// (17, 9, 'neigh_op_rgt_0')
// (17, 10, 'neigh_op_bnr_0')
// (18, 8, 'neigh_op_top_0')
// (18, 9, 'lutff_0/out')
// (18, 10, 'neigh_op_bot_0')
// (19, 8, 'neigh_op_tnl_0')
// (19, 9, 'neigh_op_lft_0')
// (19, 10, 'neigh_op_bnl_0')

reg n1156 = 0;
// (17, 8, 'local_g2_5')
// (17, 8, 'lutff_2/in_3')
// (17, 8, 'neigh_op_tnr_5')
// (17, 9, 'neigh_op_rgt_5')
// (17, 10, 'neigh_op_bnr_5')
// (18, 8, 'neigh_op_top_5')
// (18, 9, 'lutff_5/out')
// (18, 10, 'neigh_op_bot_5')
// (19, 8, 'neigh_op_tnl_5')
// (19, 9, 'neigh_op_lft_5')
// (19, 10, 'neigh_op_bnl_5')

reg n1157 = 0;
// (17, 8, 'local_g3_1')
// (17, 8, 'lutff_1/in_3')
// (17, 8, 'neigh_op_tnr_1')
// (17, 9, 'neigh_op_rgt_1')
// (17, 10, 'neigh_op_bnr_1')
// (18, 8, 'neigh_op_top_1')
// (18, 9, 'lutff_1/out')
// (18, 10, 'neigh_op_bot_1')
// (19, 8, 'neigh_op_tnl_1')
// (19, 9, 'neigh_op_lft_1')
// (19, 10, 'neigh_op_bnl_1')

reg n1158 = 0;
// (17, 8, 'local_g3_6')
// (17, 8, 'lutff_4/in_3')
// (17, 8, 'neigh_op_tnr_6')
// (17, 9, 'neigh_op_rgt_6')
// (17, 10, 'neigh_op_bnr_6')
// (18, 8, 'neigh_op_top_6')
// (18, 9, 'lutff_6/out')
// (18, 10, 'neigh_op_bot_6')
// (19, 8, 'neigh_op_tnl_6')
// (19, 9, 'neigh_op_lft_6')
// (19, 10, 'neigh_op_bnl_6')

reg n1159 = 0;
// (17, 10, 'neigh_op_tnr_0')
// (17, 11, 'neigh_op_rgt_0')
// (17, 12, 'local_g0_0')
// (17, 12, 'lutff_5/in_1')
// (17, 12, 'neigh_op_bnr_0')
// (18, 10, 'neigh_op_top_0')
// (18, 11, 'lutff_0/out')
// (18, 12, 'neigh_op_bot_0')
// (19, 10, 'neigh_op_tnl_0')
// (19, 11, 'neigh_op_lft_0')
// (19, 12, 'neigh_op_bnl_0')

reg n1160 = 0;
// (17, 10, 'neigh_op_tnr_1')
// (17, 11, 'neigh_op_rgt_1')
// (17, 12, 'local_g0_1')
// (17, 12, 'lutff_6/in_1')
// (17, 12, 'neigh_op_bnr_1')
// (18, 10, 'neigh_op_top_1')
// (18, 11, 'lutff_1/out')
// (18, 12, 'neigh_op_bot_1')
// (19, 10, 'neigh_op_tnl_1')
// (19, 11, 'neigh_op_lft_1')
// (19, 12, 'neigh_op_bnl_1')

reg n1161 = 0;
// (17, 10, 'neigh_op_tnr_2')
// (17, 11, 'neigh_op_rgt_2')
// (17, 12, 'local_g0_2')
// (17, 12, 'lutff_7/in_3')
// (17, 12, 'neigh_op_bnr_2')
// (18, 10, 'neigh_op_top_2')
// (18, 11, 'lutff_2/out')
// (18, 12, 'neigh_op_bot_2')
// (19, 10, 'neigh_op_tnl_2')
// (19, 11, 'neigh_op_lft_2')
// (19, 12, 'neigh_op_bnl_2')

reg n1162 = 0;
// (17, 10, 'neigh_op_tnr_3')
// (17, 11, 'neigh_op_rgt_3')
// (17, 12, 'neigh_op_bnr_3')
// (18, 10, 'neigh_op_top_3')
// (18, 10, 'sp12_v_t_22')
// (18, 11, 'lutff_3/out')
// (18, 11, 'sp12_v_b_22')
// (18, 12, 'neigh_op_bot_3')
// (18, 12, 'sp12_v_b_21')
// (18, 13, 'sp12_v_b_18')
// (18, 14, 'sp12_v_b_17')
// (18, 15, 'sp12_v_b_14')
// (18, 16, 'sp12_v_b_13')
// (18, 17, 'sp12_v_b_10')
// (18, 18, 'sp12_v_b_9')
// (18, 19, 'sp12_v_b_6')
// (18, 20, 'sp12_v_b_5')
// (18, 21, 'sp12_v_b_2')
// (18, 22, 'sp12_v_b_1')
// (18, 22, 'sp12_v_t_22')
// (18, 23, 'sp12_v_b_22')
// (18, 24, 'local_g2_5')
// (18, 24, 'lutff_2/in_3')
// (18, 24, 'sp12_v_b_21')
// (18, 25, 'sp12_v_b_18')
// (18, 26, 'sp12_v_b_17')
// (18, 27, 'sp12_v_b_14')
// (18, 28, 'sp12_v_b_13')
// (18, 29, 'sp12_v_b_10')
// (18, 30, 'sp12_v_b_9')
// (18, 31, 'sp12_v_b_6')
// (18, 32, 'sp12_v_b_5')
// (18, 33, 'span12_vert_2')
// (19, 10, 'neigh_op_tnl_3')
// (19, 11, 'neigh_op_lft_3')
// (19, 12, 'neigh_op_bnl_3')

reg n1163 = 0;
// (17, 10, 'sp4_h_r_10')
// (18, 9, 'neigh_op_tnr_1')
// (18, 10, 'neigh_op_rgt_1')
// (18, 10, 'sp4_h_r_23')
// (18, 11, 'neigh_op_bnr_1')
// (19, 9, 'neigh_op_top_1')
// (19, 10, 'lutff_1/out')
// (19, 10, 'sp4_h_r_34')
// (19, 11, 'neigh_op_bot_1')
// (20, 9, 'neigh_op_tnl_1')
// (20, 10, 'neigh_op_lft_1')
// (20, 10, 'sp4_h_r_47')
// (20, 11, 'neigh_op_bnl_1')
// (20, 11, 'sp4_r_v_b_47')
// (20, 12, 'sp4_r_v_b_34')
// (20, 13, 'sp4_r_v_b_23')
// (20, 14, 'sp4_r_v_b_10')
// (21, 10, 'sp4_h_l_47')
// (21, 10, 'sp4_v_t_47')
// (21, 11, 'sp4_v_b_47')
// (21, 12, 'sp4_v_b_34')
// (21, 13, 'local_g1_7')
// (21, 13, 'lutff_7/in_1')
// (21, 13, 'sp4_v_b_23')
// (21, 14, 'sp4_v_b_10')

reg n1164 = 0;
// (17, 10, 'sp4_r_v_b_40')
// (17, 11, 'sp4_r_v_b_29')
// (17, 12, 'sp4_r_v_b_16')
// (17, 13, 'sp4_r_v_b_5')
// (17, 14, 'sp4_r_v_b_40')
// (17, 15, 'sp4_r_v_b_29')
// (17, 16, 'local_g3_0')
// (17, 16, 'lutff_4/in_1')
// (17, 16, 'sp4_r_v_b_16')
// (17, 17, 'sp4_r_v_b_5')
// (18, 8, 'neigh_op_tnr_0')
// (18, 9, 'neigh_op_rgt_0')
// (18, 9, 'sp4_h_r_5')
// (18, 9, 'sp4_v_t_40')
// (18, 10, 'neigh_op_bnr_0')
// (18, 10, 'sp4_v_b_40')
// (18, 11, 'sp4_v_b_29')
// (18, 12, 'sp4_v_b_16')
// (18, 13, 'sp4_v_b_5')
// (18, 13, 'sp4_v_t_40')
// (18, 14, 'sp4_v_b_40')
// (18, 15, 'sp4_v_b_29')
// (18, 16, 'sp4_v_b_16')
// (18, 17, 'sp4_v_b_5')
// (19, 8, 'neigh_op_top_0')
// (19, 9, 'lutff_0/out')
// (19, 9, 'sp4_h_r_16')
// (19, 10, 'neigh_op_bot_0')
// (20, 8, 'neigh_op_tnl_0')
// (20, 9, 'neigh_op_lft_0')
// (20, 9, 'sp4_h_r_29')
// (20, 10, 'neigh_op_bnl_0')
// (21, 9, 'sp4_h_r_40')
// (22, 9, 'sp4_h_l_40')

reg n1165 = 0;
// (17, 10, 'sp4_r_v_b_44')
// (17, 11, 'neigh_op_tnr_2')
// (17, 11, 'sp4_r_v_b_33')
// (17, 12, 'neigh_op_rgt_2')
// (17, 12, 'sp4_r_v_b_20')
// (17, 13, 'neigh_op_bnr_2')
// (17, 13, 'sp4_r_v_b_9')
// (18, 9, 'sp4_v_t_44')
// (18, 10, 'sp4_v_b_44')
// (18, 11, 'neigh_op_top_2')
// (18, 11, 'sp4_v_b_33')
// (18, 12, 'lutff_2/out')
// (18, 12, 'sp4_v_b_20')
// (18, 13, 'neigh_op_bot_2')
// (18, 13, 'sp4_h_r_9')
// (18, 13, 'sp4_v_b_9')
// (19, 11, 'neigh_op_tnl_2')
// (19, 12, 'neigh_op_lft_2')
// (19, 13, 'neigh_op_bnl_2')
// (19, 13, 'sp4_h_r_20')
// (20, 13, 'sp4_h_r_33')
// (21, 13, 'local_g2_4')
// (21, 13, 'lutff_1/in_3')
// (21, 13, 'sp4_h_r_44')
// (22, 13, 'sp4_h_l_44')

reg n1166 = 0;
// (17, 11, 'local_g0_4')
// (17, 11, 'lutff_5/in_3')
// (17, 11, 'sp4_h_r_4')
// (18, 10, 'neigh_op_tnr_6')
// (18, 11, 'neigh_op_rgt_6')
// (18, 11, 'sp4_h_r_17')
// (18, 12, 'neigh_op_bnr_6')
// (19, 10, 'neigh_op_top_6')
// (19, 11, 'lutff_6/out')
// (19, 11, 'sp4_h_r_28')
// (19, 12, 'neigh_op_bot_6')
// (20, 10, 'neigh_op_tnl_6')
// (20, 11, 'neigh_op_lft_6')
// (20, 11, 'sp4_h_r_41')
// (20, 12, 'neigh_op_bnl_6')
// (21, 11, 'sp4_h_l_41')

reg n1167 = 0;
// (17, 11, 'local_g1_2')
// (17, 11, 'lutff_0/in_3')
// (17, 11, 'sp4_h_r_2')
// (18, 10, 'neigh_op_tnr_5')
// (18, 11, 'neigh_op_rgt_5')
// (18, 11, 'sp4_h_r_15')
// (18, 12, 'neigh_op_bnr_5')
// (19, 10, 'neigh_op_top_5')
// (19, 11, 'lutff_5/out')
// (19, 11, 'sp4_h_r_26')
// (19, 12, 'neigh_op_bot_5')
// (20, 10, 'neigh_op_tnl_5')
// (20, 11, 'neigh_op_lft_5')
// (20, 11, 'sp4_h_r_39')
// (20, 12, 'neigh_op_bnl_5')
// (21, 11, 'sp4_h_l_39')

wire n1168;
// (17, 11, 'lutff_1/lout')
// (17, 11, 'lutff_2/in_2')

wire n1169;
// (17, 11, 'lutff_3/lout')
// (17, 11, 'lutff_4/in_2')

reg n1170 = 0;
// (17, 11, 'neigh_op_tnr_0')
// (17, 12, 'neigh_op_rgt_0')
// (17, 13, 'neigh_op_bnr_0')
// (18, 8, 'sp12_v_t_23')
// (18, 9, 'sp12_v_b_23')
// (18, 10, 'sp12_v_b_20')
// (18, 11, 'neigh_op_top_0')
// (18, 11, 'sp12_v_b_19')
// (18, 12, 'lutff_0/out')
// (18, 12, 'sp12_v_b_16')
// (18, 13, 'neigh_op_bot_0')
// (18, 13, 'sp12_v_b_15')
// (18, 14, 'sp12_v_b_12')
// (18, 15, 'local_g2_3')
// (18, 15, 'lutff_4/in_3')
// (18, 15, 'sp12_v_b_11')
// (18, 16, 'sp12_v_b_8')
// (18, 17, 'sp12_v_b_7')
// (18, 18, 'sp12_v_b_4')
// (18, 19, 'sp12_v_b_3')
// (18, 20, 'sp12_v_b_0')
// (19, 11, 'neigh_op_tnl_0')
// (19, 12, 'neigh_op_lft_0')
// (19, 13, 'neigh_op_bnl_0')

reg n1171 = 0;
// (17, 11, 'neigh_op_tnr_1')
// (17, 12, 'neigh_op_rgt_1')
// (17, 13, 'neigh_op_bnr_1')
// (18, 11, 'neigh_op_top_1')
// (18, 12, 'lutff_1/out')
// (18, 13, 'neigh_op_bot_1')
// (19, 11, 'neigh_op_tnl_1')
// (19, 12, 'neigh_op_lft_1')
// (19, 13, 'local_g3_1')
// (19, 13, 'lutff_7/in_3')
// (19, 13, 'neigh_op_bnl_1')

reg n1172 = 0;
// (17, 11, 'neigh_op_tnr_3')
// (17, 12, 'neigh_op_rgt_3')
// (17, 12, 'sp4_h_r_11')
// (17, 13, 'neigh_op_bnr_3')
// (18, 11, 'neigh_op_top_3')
// (18, 12, 'lutff_3/out')
// (18, 12, 'sp4_h_r_22')
// (18, 13, 'neigh_op_bot_3')
// (19, 11, 'neigh_op_tnl_3')
// (19, 12, 'neigh_op_lft_3')
// (19, 12, 'sp4_h_r_35')
// (19, 13, 'neigh_op_bnl_3')
// (20, 12, 'sp4_h_r_46')
// (20, 13, 'sp4_r_v_b_46')
// (20, 14, 'sp4_r_v_b_35')
// (20, 15, 'sp4_r_v_b_22')
// (20, 16, 'sp4_r_v_b_11')
// (21, 12, 'sp4_h_l_46')
// (21, 12, 'sp4_v_t_46')
// (21, 13, 'sp4_v_b_46')
// (21, 14, 'sp4_v_b_35')
// (21, 15, 'sp4_v_b_22')
// (21, 16, 'local_g0_3')
// (21, 16, 'lutff_5/in_2')
// (21, 16, 'sp4_v_b_11')

reg n1173 = 0;
// (17, 11, 'neigh_op_tnr_4')
// (17, 12, 'neigh_op_rgt_4')
// (17, 13, 'neigh_op_bnr_4')
// (18, 11, 'neigh_op_top_4')
// (18, 12, 'lutff_4/out')
// (18, 12, 'sp4_h_r_8')
// (18, 13, 'neigh_op_bot_4')
// (19, 11, 'neigh_op_tnl_4')
// (19, 12, 'neigh_op_lft_4')
// (19, 12, 'sp4_h_r_21')
// (19, 13, 'neigh_op_bnl_4')
// (20, 12, 'sp4_h_r_32')
// (21, 12, 'sp4_h_r_45')
// (21, 13, 'sp4_r_v_b_36')
// (21, 14, 'sp4_r_v_b_25')
// (21, 15, 'sp4_r_v_b_12')
// (21, 16, 'sp4_r_v_b_1')
// (22, 12, 'sp4_h_l_45')
// (22, 12, 'sp4_v_t_36')
// (22, 13, 'sp4_v_b_36')
// (22, 14, 'sp4_v_b_25')
// (22, 15, 'sp4_v_b_12')
// (22, 16, 'local_g1_1')
// (22, 16, 'lutff_3/in_3')
// (22, 16, 'sp4_v_b_1')

reg n1174 = 0;
// (17, 11, 'neigh_op_tnr_5')
// (17, 12, 'neigh_op_rgt_5')
// (17, 13, 'neigh_op_bnr_5')
// (18, 11, 'neigh_op_top_5')
// (18, 12, 'lutff_5/out')
// (18, 12, 'sp4_r_v_b_43')
// (18, 13, 'neigh_op_bot_5')
// (18, 13, 'sp4_r_v_b_30')
// (18, 14, 'sp4_r_v_b_19')
// (18, 15, 'sp4_r_v_b_6')
// (18, 16, 'sp4_r_v_b_39')
// (18, 17, 'sp4_r_v_b_26')
// (18, 18, 'sp4_r_v_b_15')
// (18, 19, 'sp4_r_v_b_2')
// (19, 11, 'neigh_op_tnl_5')
// (19, 11, 'sp4_v_t_43')
// (19, 12, 'neigh_op_lft_5')
// (19, 12, 'sp4_v_b_43')
// (19, 13, 'neigh_op_bnl_5')
// (19, 13, 'sp4_v_b_30')
// (19, 14, 'sp4_v_b_19')
// (19, 15, 'sp4_v_b_6')
// (19, 15, 'sp4_v_t_39')
// (19, 16, 'sp4_v_b_39')
// (19, 17, 'sp4_v_b_26')
// (19, 18, 'local_g1_7')
// (19, 18, 'lutff_7/in_3')
// (19, 18, 'sp4_v_b_15')
// (19, 19, 'sp4_v_b_2')

reg n1175 = 0;
// (17, 11, 'neigh_op_tnr_6')
// (17, 12, 'neigh_op_rgt_6')
// (17, 13, 'neigh_op_bnr_6')
// (18, 11, 'neigh_op_top_6')
// (18, 12, 'lutff_6/out')
// (18, 12, 'sp4_r_v_b_45')
// (18, 13, 'neigh_op_bot_6')
// (18, 13, 'sp4_r_v_b_32')
// (18, 14, 'sp4_r_v_b_21')
// (18, 15, 'sp4_r_v_b_8')
// (19, 11, 'neigh_op_tnl_6')
// (19, 11, 'sp4_v_t_45')
// (19, 12, 'neigh_op_lft_6')
// (19, 12, 'sp4_v_b_45')
// (19, 13, 'neigh_op_bnl_6')
// (19, 13, 'sp4_v_b_32')
// (19, 14, 'local_g1_5')
// (19, 14, 'lutff_7/in_3')
// (19, 14, 'sp4_v_b_21')
// (19, 15, 'sp4_v_b_8')

reg n1176 = 0;
// (17, 11, 'neigh_op_tnr_7')
// (17, 12, 'neigh_op_rgt_7')
// (17, 13, 'local_g1_7')
// (17, 13, 'lutff_6/in_0')
// (17, 13, 'neigh_op_bnr_7')
// (18, 11, 'neigh_op_top_7')
// (18, 12, 'lutff_7/out')
// (18, 13, 'neigh_op_bot_7')
// (19, 11, 'neigh_op_tnl_7')
// (19, 12, 'neigh_op_lft_7')
// (19, 13, 'neigh_op_bnl_7')

reg n1177 = 0;
// (17, 11, 'sp12_h_r_0')
// (17, 11, 'sp12_v_t_23')
// (17, 12, 'sp12_v_b_23')
// (17, 13, 'sp12_v_b_20')
// (17, 14, 'sp12_v_b_19')
// (17, 15, 'sp12_v_b_16')
// (17, 16, 'sp12_v_b_15')
// (17, 17, 'local_g2_4')
// (17, 17, 'lutff_1/in_1')
// (17, 17, 'sp12_v_b_12')
// (17, 18, 'sp12_v_b_11')
// (17, 19, 'sp12_v_b_8')
// (17, 20, 'sp12_v_b_7')
// (17, 21, 'sp12_v_b_4')
// (17, 22, 'sp12_v_b_3')
// (17, 23, 'sp12_v_b_0')
// (18, 11, 'sp12_h_r_3')
// (19, 11, 'sp12_h_r_4')
// (20, 10, 'neigh_op_tnr_0')
// (20, 11, 'neigh_op_rgt_0')
// (20, 11, 'sp12_h_r_7')
// (20, 12, 'neigh_op_bnr_0')
// (21, 10, 'neigh_op_top_0')
// (21, 11, 'lutff_0/out')
// (21, 11, 'sp12_h_r_8')
// (21, 12, 'neigh_op_bot_0')
// (22, 10, 'neigh_op_tnl_0')
// (22, 11, 'neigh_op_lft_0')
// (22, 11, 'sp12_h_r_11')
// (22, 12, 'neigh_op_bnl_0')
// (23, 11, 'sp12_h_r_12')
// (24, 11, 'sp12_h_r_15')
// (25, 11, 'sp12_h_r_16')
// (26, 11, 'sp12_h_r_19')
// (27, 11, 'sp12_h_r_20')
// (28, 11, 'sp12_h_r_23')
// (29, 11, 'sp12_h_l_23')

reg n1178 = 0;
// (17, 11, 'sp4_h_r_0')
// (18, 10, 'neigh_op_tnr_4')
// (18, 11, 'neigh_op_rgt_4')
// (18, 11, 'sp4_h_r_13')
// (18, 12, 'neigh_op_bnr_4')
// (19, 10, 'neigh_op_top_4')
// (19, 11, 'lutff_4/out')
// (19, 11, 'sp4_h_r_24')
// (19, 12, 'neigh_op_bot_4')
// (20, 10, 'neigh_op_tnl_4')
// (20, 11, 'neigh_op_lft_4')
// (20, 11, 'sp4_h_r_37')
// (20, 12, 'neigh_op_bnl_4')
// (20, 12, 'sp4_r_v_b_37')
// (20, 13, 'sp4_r_v_b_24')
// (20, 14, 'sp4_r_v_b_13')
// (20, 15, 'sp4_r_v_b_0')
// (21, 11, 'sp4_h_l_37')
// (21, 11, 'sp4_v_t_37')
// (21, 12, 'sp4_v_b_37')
// (21, 13, 'sp4_v_b_24')
// (21, 14, 'sp4_v_b_13')
// (21, 15, 'local_g1_0')
// (21, 15, 'lutff_6/in_3')
// (21, 15, 'sp4_v_b_0')

wire n1179;
// (17, 11, 'sp4_h_r_7')
// (17, 15, 'sp4_h_r_3')
// (18, 11, 'local_g0_2')
// (18, 11, 'lutff_global/cen')
// (18, 11, 'sp4_h_r_18')
// (18, 15, 'sp4_h_r_14')
// (19, 11, 'sp4_h_r_31')
// (19, 14, 'neigh_op_tnr_3')
// (19, 15, 'neigh_op_rgt_3')
// (19, 15, 'sp4_h_r_27')
// (19, 16, 'neigh_op_bnr_3')
// (20, 11, 'sp4_h_r_42')
// (20, 12, 'sp4_r_v_b_42')
// (20, 13, 'sp4_r_v_b_31')
// (20, 14, 'neigh_op_top_3')
// (20, 14, 'sp4_r_v_b_18')
// (20, 15, 'lutff_3/out')
// (20, 15, 'sp4_h_r_38')
// (20, 15, 'sp4_r_v_b_7')
// (20, 16, 'neigh_op_bot_3')
// (20, 16, 'sp4_r_v_b_38')
// (20, 17, 'sp4_r_v_b_27')
// (20, 18, 'sp4_r_v_b_14')
// (20, 19, 'sp4_r_v_b_3')
// (21, 11, 'sp4_h_l_42')
// (21, 11, 'sp4_v_t_42')
// (21, 12, 'sp4_v_b_42')
// (21, 13, 'sp4_v_b_31')
// (21, 14, 'neigh_op_tnl_3')
// (21, 14, 'sp4_v_b_18')
// (21, 15, 'neigh_op_lft_3')
// (21, 15, 'sp4_h_l_38')
// (21, 15, 'sp4_v_b_7')
// (21, 15, 'sp4_v_t_38')
// (21, 16, 'neigh_op_bnl_3')
// (21, 16, 'sp4_v_b_38')
// (21, 17, 'local_g3_3')
// (21, 17, 'lutff_global/cen')
// (21, 17, 'sp4_v_b_27')
// (21, 18, 'sp4_v_b_14')
// (21, 19, 'sp4_v_b_3')

reg n1180 = 0;
// (17, 11, 'sp4_r_v_b_37')
// (17, 11, 'sp4_r_v_b_45')
// (17, 12, 'local_g0_3')
// (17, 12, 'lutff_1/in_0')
// (17, 12, 'sp4_r_v_b_24')
// (17, 12, 'sp4_r_v_b_32')
// (17, 13, 'local_g2_5')
// (17, 13, 'lutff_1/in_0')
// (17, 13, 'lutff_5/in_0')
// (17, 13, 'lutff_6/in_1')
// (17, 13, 'sp4_r_v_b_13')
// (17, 13, 'sp4_r_v_b_21')
// (17, 14, 'local_g1_0')
// (17, 14, 'local_g2_0')
// (17, 14, 'lutff_0/in_0')
// (17, 14, 'lutff_3/in_0')
// (17, 14, 'lutff_6/in_0')
// (17, 14, 'sp4_r_v_b_0')
// (17, 14, 'sp4_r_v_b_8')
// (17, 15, 'local_g2_4')
// (17, 15, 'local_g3_4')
// (17, 15, 'lutff_0/in_0')
// (17, 15, 'lutff_3/in_0')
// (17, 15, 'lutff_5/in_0')
// (17, 15, 'lutff_7/in_0')
// (17, 15, 'neigh_op_tnr_4')
// (17, 15, 'sp4_r_v_b_37')
// (17, 16, 'local_g0_0')
// (17, 16, 'local_g3_4')
// (17, 16, 'lutff_1/in_0')
// (17, 16, 'lutff_2/in_0')
// (17, 16, 'neigh_op_rgt_4')
// (17, 16, 'sp4_r_v_b_24')
// (17, 17, 'local_g0_4')
// (17, 17, 'lutff_6/in_0')
// (17, 17, 'neigh_op_bnr_4')
// (17, 17, 'sp4_r_v_b_13')
// (17, 18, 'sp4_r_v_b_0')
// (18, 10, 'sp4_v_t_37')
// (18, 10, 'sp4_v_t_45')
// (18, 11, 'sp4_v_b_37')
// (18, 11, 'sp4_v_b_45')
// (18, 12, 'sp4_r_v_b_37')
// (18, 12, 'sp4_v_b_24')
// (18, 12, 'sp4_v_b_32')
// (18, 13, 'sp4_r_v_b_24')
// (18, 13, 'sp4_v_b_13')
// (18, 13, 'sp4_v_b_21')
// (18, 14, 'sp4_h_r_5')
// (18, 14, 'sp4_r_v_b_13')
// (18, 14, 'sp4_v_b_0')
// (18, 14, 'sp4_v_b_8')
// (18, 14, 'sp4_v_t_37')
// (18, 15, 'local_g2_4')
// (18, 15, 'lutff_2/in_0')
// (18, 15, 'lutff_4/in_2')
// (18, 15, 'neigh_op_top_4')
// (18, 15, 'sp4_r_v_b_0')
// (18, 15, 'sp4_r_v_b_36')
// (18, 15, 'sp4_v_b_37')
// (18, 16, 'local_g0_4')
// (18, 16, 'lutff_4/in_0')
// (18, 16, 'lutff_4/out')
// (18, 16, 'sp4_r_v_b_25')
// (18, 16, 'sp4_r_v_b_41')
// (18, 16, 'sp4_v_b_24')
// (18, 17, 'neigh_op_bot_4')
// (18, 17, 'sp4_r_v_b_12')
// (18, 17, 'sp4_r_v_b_28')
// (18, 17, 'sp4_v_b_13')
// (18, 18, 'sp4_r_v_b_1')
// (18, 18, 'sp4_r_v_b_17')
// (18, 18, 'sp4_v_b_0')
// (18, 19, 'sp4_r_v_b_4')
// (19, 11, 'sp4_v_t_37')
// (19, 12, 'sp4_v_b_37')
// (19, 13, 'local_g3_0')
// (19, 13, 'lutff_1/in_2')
// (19, 13, 'lutff_5/in_0')
// (19, 13, 'lutff_7/in_0')
// (19, 13, 'sp4_v_b_24')
// (19, 14, 'local_g0_5')
// (19, 14, 'lutff_1/in_0')
// (19, 14, 'lutff_3/in_2')
// (19, 14, 'lutff_7/in_0')
// (19, 14, 'sp4_h_r_16')
// (19, 14, 'sp4_v_b_13')
// (19, 14, 'sp4_v_t_36')
// (19, 15, 'local_g2_4')
// (19, 15, 'local_g3_4')
// (19, 15, 'lutff_1/in_0')
// (19, 15, 'lutff_3/in_0')
// (19, 15, 'lutff_6/in_0')
// (19, 15, 'neigh_op_tnl_4')
// (19, 15, 'sp4_v_b_0')
// (19, 15, 'sp4_v_b_36')
// (19, 15, 'sp4_v_t_41')
// (19, 16, 'neigh_op_lft_4')
// (19, 16, 'sp4_v_b_25')
// (19, 16, 'sp4_v_b_41')
// (19, 17, 'neigh_op_bnl_4')
// (19, 17, 'sp4_v_b_12')
// (19, 17, 'sp4_v_b_28')
// (19, 18, 'local_g0_1')
// (19, 18, 'lutff_1/in_0')
// (19, 18, 'lutff_3/in_0')
// (19, 18, 'lutff_7/in_0')
// (19, 18, 'sp4_h_r_1')
// (19, 18, 'sp4_v_b_1')
// (19, 18, 'sp4_v_b_17')
// (19, 19, 'sp4_h_r_4')
// (19, 19, 'sp4_v_b_4')
// (20, 14, 'sp4_h_r_29')
// (20, 18, 'sp4_h_r_12')
// (20, 19, 'sp4_h_r_17')
// (21, 11, 'sp4_r_v_b_40')
// (21, 12, 'sp4_r_v_b_29')
// (21, 13, 'local_g3_0')
// (21, 13, 'lutff_1/in_0')
// (21, 13, 'lutff_5/in_0')
// (21, 13, 'lutff_7/in_0')
// (21, 13, 'sp4_r_v_b_16')
// (21, 14, 'local_g3_0')
// (21, 14, 'lutff_0/in_1')
// (21, 14, 'lutff_3/in_0')
// (21, 14, 'lutff_6/in_1')
// (21, 14, 'sp4_h_r_40')
// (21, 14, 'sp4_r_v_b_5')
// (21, 15, 'sp4_r_v_b_40')
// (21, 16, 'local_g0_5')
// (21, 16, 'lutff_1/in_0')
// (21, 16, 'lutff_3/in_0')
// (21, 16, 'lutff_5/in_0')
// (21, 16, 'sp4_r_v_b_29')
// (21, 17, 'sp4_r_v_b_16')
// (21, 18, 'local_g2_1')
// (21, 18, 'local_g3_1')
// (21, 18, 'lutff_0/in_0')
// (21, 18, 'lutff_3/in_0')
// (21, 18, 'lutff_6/in_0')
// (21, 18, 'sp4_h_r_25')
// (21, 18, 'sp4_r_v_b_5')
// (21, 19, 'sp4_h_r_28')
// (22, 10, 'sp4_v_t_40')
// (22, 11, 'sp4_v_b_40')
// (22, 12, 'sp4_v_b_29')
// (22, 13, 'local_g0_0')
// (22, 13, 'local_g1_0')
// (22, 13, 'lutff_0/in_0')
// (22, 13, 'lutff_3/in_0')
// (22, 13, 'lutff_6/in_0')
// (22, 13, 'sp4_v_b_16')
// (22, 14, 'sp4_h_l_40')
// (22, 14, 'sp4_v_b_5')
// (22, 14, 'sp4_v_t_40')
// (22, 15, 'sp4_v_b_40')
// (22, 16, 'local_g2_5')
// (22, 16, 'lutff_1/in_0')
// (22, 16, 'lutff_3/in_0')
// (22, 16, 'lutff_5/in_0')
// (22, 16, 'sp4_r_v_b_41')
// (22, 16, 'sp4_r_v_b_47')
// (22, 16, 'sp4_v_b_29')
// (22, 17, 'sp4_r_v_b_28')
// (22, 17, 'sp4_r_v_b_34')
// (22, 17, 'sp4_v_b_16')
// (22, 18, 'sp4_h_r_36')
// (22, 18, 'sp4_r_v_b_17')
// (22, 18, 'sp4_r_v_b_23')
// (22, 18, 'sp4_v_b_5')
// (22, 19, 'sp4_h_r_41')
// (22, 19, 'sp4_r_v_b_10')
// (22, 19, 'sp4_r_v_b_4')
// (23, 15, 'sp4_v_t_41')
// (23, 15, 'sp4_v_t_47')
// (23, 16, 'sp4_v_b_41')
// (23, 16, 'sp4_v_b_47')
// (23, 17, 'local_g2_4')
// (23, 17, 'local_g3_2')
// (23, 17, 'lutff_1/in_0')
// (23, 17, 'lutff_3/in_0')
// (23, 17, 'lutff_6/in_0')
// (23, 17, 'sp4_v_b_28')
// (23, 17, 'sp4_v_b_34')
// (23, 18, 'sp4_h_l_36')
// (23, 18, 'sp4_v_b_17')
// (23, 18, 'sp4_v_b_23')
// (23, 19, 'sp4_h_l_41')
// (23, 19, 'sp4_v_b_10')
// (23, 19, 'sp4_v_b_4')

reg n1181 = 0;
// (17, 12, 'local_g1_3')
// (17, 12, 'lutff_3/in_1')
// (17, 12, 'sp4_h_r_3')
// (18, 12, 'sp4_h_r_14')
// (19, 12, 'sp4_h_r_27')
// (20, 9, 'sp4_r_v_b_38')
// (20, 10, 'neigh_op_tnr_7')
// (20, 10, 'sp4_r_v_b_27')
// (20, 11, 'neigh_op_rgt_7')
// (20, 11, 'sp4_r_v_b_14')
// (20, 12, 'neigh_op_bnr_7')
// (20, 12, 'sp4_h_r_38')
// (20, 12, 'sp4_r_v_b_3')
// (21, 8, 'sp4_v_t_38')
// (21, 9, 'sp4_v_b_38')
// (21, 10, 'neigh_op_top_7')
// (21, 10, 'sp4_v_b_27')
// (21, 11, 'lutff_7/out')
// (21, 11, 'sp4_v_b_14')
// (21, 12, 'neigh_op_bot_7')
// (21, 12, 'sp4_h_l_38')
// (21, 12, 'sp4_v_b_3')
// (22, 10, 'neigh_op_tnl_7')
// (22, 11, 'neigh_op_lft_7')
// (22, 12, 'neigh_op_bnl_7')

wire n1182;
// (17, 12, 'lutff_1/lout')
// (17, 12, 'lutff_2/in_2')

wire n1183;
// (17, 12, 'neigh_op_tnr_4')
// (17, 13, 'neigh_op_rgt_4')
// (17, 14, 'neigh_op_bnr_4')
// (18, 12, 'neigh_op_top_4')
// (18, 13, 'local_g1_4')
// (18, 13, 'lutff_0/in_1')
// (18, 13, 'lutff_4/out')
// (18, 14, 'neigh_op_bot_4')
// (19, 12, 'neigh_op_tnl_4')
// (19, 13, 'neigh_op_lft_4')
// (19, 14, 'neigh_op_bnl_4')

wire n1184;
// (17, 12, 'neigh_op_tnr_7')
// (17, 13, 'neigh_op_rgt_7')
// (17, 14, 'neigh_op_bnr_7')
// (18, 12, 'neigh_op_top_7')
// (18, 13, 'local_g2_7')
// (18, 13, 'lutff_0/in_3')
// (18, 13, 'lutff_7/out')
// (18, 14, 'neigh_op_bot_7')
// (19, 12, 'neigh_op_tnl_7')
// (19, 13, 'neigh_op_lft_7')
// (19, 14, 'neigh_op_bnl_7')

reg n1185 = 0;
// (17, 12, 'sp4_h_r_1')
// (18, 12, 'sp4_h_r_12')
// (19, 11, 'neigh_op_tnr_2')
// (19, 12, 'neigh_op_rgt_2')
// (19, 12, 'sp4_h_r_25')
// (19, 13, 'neigh_op_bnr_2')
// (20, 11, 'neigh_op_top_2')
// (20, 12, 'lutff_2/out')
// (20, 12, 'sp4_h_r_36')
// (20, 13, 'neigh_op_bot_2')
// (20, 13, 'sp4_r_v_b_36')
// (20, 14, 'sp4_r_v_b_25')
// (20, 15, 'sp4_r_v_b_12')
// (20, 16, 'sp4_r_v_b_1')
// (21, 11, 'neigh_op_tnl_2')
// (21, 12, 'neigh_op_lft_2')
// (21, 12, 'sp4_h_l_36')
// (21, 12, 'sp4_v_t_36')
// (21, 13, 'neigh_op_bnl_2')
// (21, 13, 'sp4_v_b_36')
// (21, 14, 'local_g3_1')
// (21, 14, 'lutff_7/in_3')
// (21, 14, 'sp4_v_b_25')
// (21, 15, 'sp4_v_b_12')
// (21, 16, 'sp4_v_b_1')

wire n1186;
// (17, 12, 'sp4_h_r_8')
// (18, 11, 'neigh_op_tnr_0')
// (18, 12, 'neigh_op_rgt_0')
// (18, 12, 'sp4_h_r_21')
// (18, 13, 'neigh_op_bnr_0')
// (19, 11, 'neigh_op_top_0')
// (19, 12, 'lutff_0/out')
// (19, 12, 'sp4_h_r_32')
// (19, 13, 'neigh_op_bot_0')
// (20, 11, 'neigh_op_tnl_0')
// (20, 12, 'neigh_op_lft_0')
// (20, 12, 'sp4_h_r_45')
// (20, 13, 'neigh_op_bnl_0')
// (21, 12, 'local_g1_3')
// (21, 12, 'lutff_global/cen')
// (21, 12, 'sp4_h_l_45')
// (21, 12, 'sp4_h_r_11')
// (22, 12, 'sp4_h_r_22')
// (23, 12, 'sp4_h_r_35')
// (24, 12, 'sp4_h_r_46')
// (25, 12, 'sp4_h_l_46')

wire n1187;
// (17, 13, 'lutff_1/lout')
// (17, 13, 'lutff_2/in_2')

wire n1188;
// (17, 13, 'lutff_3/lout')
// (17, 13, 'lutff_4/in_2')

wire n1189;
// (17, 13, 'lutff_6/lout')
// (17, 13, 'lutff_7/in_2')

wire n1190;
// (17, 13, 'neigh_op_tnr_1')
// (17, 14, 'neigh_op_rgt_1')
// (17, 15, 'neigh_op_bnr_1')
// (18, 13, 'neigh_op_top_1')
// (18, 14, 'local_g2_1')
// (18, 14, 'lutff_1/out')
// (18, 14, 'lutff_6/in_1')
// (18, 15, 'neigh_op_bot_1')
// (19, 13, 'neigh_op_tnl_1')
// (19, 14, 'neigh_op_lft_1')
// (19, 15, 'neigh_op_bnl_1')

wire n1191;
// (17, 13, 'neigh_op_tnr_3')
// (17, 14, 'neigh_op_rgt_3')
// (17, 15, 'neigh_op_bnr_3')
// (18, 13, 'neigh_op_top_3')
// (18, 14, 'local_g1_3')
// (18, 14, 'lutff_1/in_3')
// (18, 14, 'lutff_3/out')
// (18, 15, 'neigh_op_bot_3')
// (19, 13, 'neigh_op_tnl_3')
// (19, 14, 'neigh_op_lft_3')
// (19, 15, 'neigh_op_bnl_3')

wire n1192;
// (17, 13, 'neigh_op_tnr_5')
// (17, 14, 'neigh_op_rgt_5')
// (17, 15, 'neigh_op_bnr_5')
// (18, 13, 'neigh_op_top_5')
// (18, 14, 'local_g2_5')
// (18, 14, 'lutff_0/in_3')
// (18, 14, 'lutff_5/out')
// (18, 15, 'neigh_op_bot_5')
// (19, 13, 'neigh_op_tnl_5')
// (19, 14, 'neigh_op_lft_5')
// (19, 15, 'neigh_op_bnl_5')

reg n1193 = 0;
// (17, 13, 'sp4_r_v_b_37')
// (17, 14, 'sp4_r_v_b_24')
// (17, 15, 'sp4_r_v_b_13')
// (17, 16, 'local_g1_0')
// (17, 16, 'lutff_3/in_0')
// (17, 16, 'sp4_r_v_b_0')
// (18, 12, 'sp4_h_r_6')
// (18, 12, 'sp4_v_t_37')
// (18, 13, 'sp4_v_b_37')
// (18, 14, 'sp4_v_b_24')
// (18, 15, 'sp4_v_b_13')
// (18, 16, 'sp4_v_b_0')
// (19, 11, 'neigh_op_tnr_7')
// (19, 12, 'neigh_op_rgt_7')
// (19, 12, 'sp4_h_r_19')
// (19, 13, 'neigh_op_bnr_7')
// (20, 11, 'neigh_op_top_7')
// (20, 12, 'lutff_7/out')
// (20, 12, 'sp4_h_r_30')
// (20, 13, 'neigh_op_bot_7')
// (21, 11, 'neigh_op_tnl_7')
// (21, 12, 'neigh_op_lft_7')
// (21, 12, 'sp4_h_r_43')
// (21, 13, 'neigh_op_bnl_7')
// (22, 12, 'sp4_h_l_43')

reg n1194 = 0;
// (17, 13, 'sp4_r_v_b_40')
// (17, 14, 'sp4_r_v_b_29')
// (17, 15, 'sp4_r_v_b_16')
// (17, 16, 'local_g1_5')
// (17, 16, 'lutff_3/in_3')
// (17, 16, 'sp4_r_v_b_5')
// (18, 12, 'sp4_h_r_11')
// (18, 12, 'sp4_v_t_40')
// (18, 13, 'sp4_v_b_40')
// (18, 14, 'sp4_v_b_29')
// (18, 15, 'sp4_v_b_16')
// (18, 16, 'sp4_v_b_5')
// (19, 12, 'sp4_h_r_22')
// (20, 11, 'neigh_op_tnr_7')
// (20, 12, 'neigh_op_rgt_7')
// (20, 12, 'sp4_h_r_35')
// (20, 13, 'neigh_op_bnr_7')
// (21, 11, 'neigh_op_top_7')
// (21, 12, 'lutff_7/out')
// (21, 12, 'sp4_h_r_46')
// (21, 13, 'neigh_op_bot_7')
// (22, 11, 'neigh_op_tnl_7')
// (22, 12, 'neigh_op_lft_7')
// (22, 12, 'sp4_h_l_46')
// (22, 13, 'neigh_op_bnl_7')

wire n1195;
// (17, 13, 'sp4_r_v_b_43')
// (17, 14, 'sp4_r_v_b_30')
// (17, 15, 'sp4_r_v_b_19')
// (17, 16, 'sp4_r_v_b_6')
// (17, 17, 'neigh_op_tnr_7')
// (17, 17, 'sp4_r_v_b_43')
// (17, 18, 'neigh_op_rgt_7')
// (17, 18, 'sp4_r_v_b_30')
// (17, 19, 'neigh_op_bnr_7')
// (17, 19, 'sp4_r_v_b_19')
// (17, 20, 'sp4_r_v_b_6')
// (18, 12, 'sp4_v_t_43')
// (18, 13, 'local_g2_3')
// (18, 13, 'lutff_4/in_3')
// (18, 13, 'sp4_v_b_43')
// (18, 14, 'sp4_v_b_30')
// (18, 15, 'sp4_v_b_19')
// (18, 16, 'sp4_v_b_6')
// (18, 16, 'sp4_v_t_43')
// (18, 17, 'neigh_op_top_7')
// (18, 17, 'sp4_v_b_43')
// (18, 18, 'lutff_7/out')
// (18, 18, 'sp4_v_b_30')
// (18, 19, 'neigh_op_bot_7')
// (18, 19, 'sp4_v_b_19')
// (18, 20, 'sp4_v_b_6')
// (19, 17, 'neigh_op_tnl_7')
// (19, 18, 'neigh_op_lft_7')
// (19, 19, 'neigh_op_bnl_7')

wire n1196;
// (17, 14, 'lutff_0/lout')
// (17, 14, 'lutff_1/in_2')

wire n1197;
// (17, 14, 'lutff_3/lout')
// (17, 14, 'lutff_4/in_2')

wire n1198;
// (17, 14, 'lutff_6/lout')
// (17, 14, 'lutff_7/in_2')

wire n1199;
// (17, 14, 'neigh_op_tnr_0')
// (17, 14, 'sp4_r_v_b_39')
// (17, 14, 'sp4_r_v_b_45')
// (17, 15, 'neigh_op_rgt_0')
// (17, 15, 'sp4_r_v_b_26')
// (17, 15, 'sp4_r_v_b_32')
// (17, 16, 'neigh_op_bnr_0')
// (17, 16, 'sp4_r_v_b_15')
// (17, 16, 'sp4_r_v_b_21')
// (17, 17, 'sp4_r_v_b_2')
// (17, 17, 'sp4_r_v_b_8')
// (18, 12, 'sp4_r_v_b_36')
// (18, 13, 'sp4_r_v_b_25')
// (18, 13, 'sp4_v_t_39')
// (18, 13, 'sp4_v_t_45')
// (18, 14, 'neigh_op_top_0')
// (18, 14, 'sp4_r_v_b_12')
// (18, 14, 'sp4_v_b_39')
// (18, 14, 'sp4_v_b_45')
// (18, 15, 'local_g2_2')
// (18, 15, 'lutff_0/out')
// (18, 15, 'lutff_global/cen')
// (18, 15, 'sp4_r_v_b_1')
// (18, 15, 'sp4_v_b_26')
// (18, 15, 'sp4_v_b_32')
// (18, 16, 'neigh_op_bot_0')
// (18, 16, 'sp4_v_b_15')
// (18, 16, 'sp4_v_b_21')
// (18, 17, 'sp4_h_r_2')
// (18, 17, 'sp4_v_b_2')
// (18, 17, 'sp4_v_b_8')
// (19, 11, 'sp4_h_r_6')
// (19, 11, 'sp4_v_t_36')
// (19, 12, 'sp4_v_b_36')
// (19, 13, 'sp4_v_b_25')
// (19, 14, 'neigh_op_tnl_0')
// (19, 14, 'sp4_v_b_12')
// (19, 15, 'neigh_op_lft_0')
// (19, 15, 'sp4_v_b_1')
// (19, 16, 'neigh_op_bnl_0')
// (19, 17, 'sp4_h_r_15')
// (20, 11, 'local_g1_3')
// (20, 11, 'lutff_global/cen')
// (20, 11, 'sp4_h_r_19')
// (20, 17, 'sp4_h_r_26')
// (21, 11, 'sp4_h_r_30')
// (21, 17, 'sp4_h_r_39')
// (22, 11, 'sp4_h_r_43')
// (22, 17, 'sp4_h_l_39')
// (23, 11, 'sp4_h_l_43')

reg n1200 = 0;
// (17, 14, 'neigh_op_tnr_1')
// (17, 15, 'neigh_op_rgt_1')
// (17, 16, 'neigh_op_bnr_1')
// (18, 14, 'neigh_op_top_1')
// (18, 15, 'local_g2_1')
// (18, 15, 'lutff_1/out')
// (18, 15, 'lutff_2/in_1')
// (18, 16, 'neigh_op_bot_1')
// (19, 14, 'neigh_op_tnl_1')
// (19, 15, 'neigh_op_lft_1')
// (19, 16, 'neigh_op_bnl_1')

wire n1201;
// (17, 14, 'neigh_op_tnr_3')
// (17, 15, 'neigh_op_rgt_3')
// (17, 16, 'neigh_op_bnr_3')
// (18, 14, 'neigh_op_top_3')
// (18, 15, 'local_g0_3')
// (18, 15, 'lutff_3/out')
// (18, 15, 'lutff_6/in_3')
// (18, 16, 'neigh_op_bot_3')
// (19, 14, 'neigh_op_tnl_3')
// (19, 15, 'neigh_op_lft_3')
// (19, 16, 'neigh_op_bnl_3')

wire n1202;
// (17, 14, 'neigh_op_tnr_6')
// (17, 15, 'neigh_op_rgt_6')
// (17, 16, 'neigh_op_bnr_6')
// (18, 14, 'local_g0_6')
// (18, 14, 'lutff_1/in_1')
// (18, 14, 'neigh_op_top_6')
// (18, 15, 'lutff_6/out')
// (18, 16, 'neigh_op_bot_6')
// (19, 14, 'neigh_op_tnl_6')
// (19, 15, 'neigh_op_lft_6')
// (19, 16, 'neigh_op_bnl_6')

reg n1203 = 0;
// (17, 15, 'local_g0_2')
// (17, 15, 'lutff_1/in_1')
// (17, 15, 'sp4_h_r_2')
// (18, 15, 'sp4_h_r_15')
// (19, 15, 'sp4_h_r_26')
// (20, 11, 'neigh_op_tnr_6')
// (20, 12, 'neigh_op_rgt_6')
// (20, 12, 'sp4_r_v_b_44')
// (20, 13, 'neigh_op_bnr_6')
// (20, 13, 'sp4_r_v_b_33')
// (20, 14, 'sp4_r_v_b_20')
// (20, 15, 'sp4_h_r_39')
// (20, 15, 'sp4_r_v_b_9')
// (21, 11, 'neigh_op_top_6')
// (21, 11, 'sp4_v_t_44')
// (21, 12, 'lutff_6/out')
// (21, 12, 'sp4_v_b_44')
// (21, 13, 'neigh_op_bot_6')
// (21, 13, 'sp4_v_b_33')
// (21, 14, 'sp4_v_b_20')
// (21, 15, 'sp4_h_l_39')
// (21, 15, 'sp4_v_b_9')
// (22, 11, 'neigh_op_tnl_6')
// (22, 12, 'neigh_op_lft_6')
// (22, 13, 'neigh_op_bnl_6')

reg n1204 = 0;
// (17, 15, 'local_g1_1')
// (17, 15, 'lutff_3/in_3')
// (17, 15, 'sp12_h_r_1')
// (18, 15, 'sp12_h_r_2')
// (19, 15, 'sp12_h_r_5')
// (20, 15, 'sp12_h_r_6')
// (21, 15, 'sp12_h_r_9')
// (22, 15, 'sp12_h_r_10')
// (23, 14, 'neigh_op_tnr_3')
// (23, 15, 'neigh_op_rgt_3')
// (23, 15, 'sp12_h_r_13')
// (23, 16, 'neigh_op_bnr_3')
// (24, 14, 'neigh_op_top_3')
// (24, 15, 'lutff_3/out')
// (24, 15, 'sp12_h_r_14')
// (24, 16, 'neigh_op_bot_3')
// (25, 14, 'neigh_op_tnl_3')
// (25, 15, 'neigh_op_lft_3')
// (25, 15, 'sp12_h_r_17')
// (25, 16, 'neigh_op_bnl_3')
// (26, 15, 'sp12_h_r_18')
// (27, 15, 'sp12_h_r_21')
// (28, 15, 'sp12_h_r_22')
// (29, 15, 'sp12_h_l_22')

wire n1205;
// (17, 15, 'lutff_0/lout')
// (17, 15, 'lutff_1/in_2')

wire n1206;
// (17, 15, 'lutff_3/lout')
// (17, 15, 'lutff_4/in_2')

wire n1207;
// (17, 15, 'lutff_5/lout')
// (17, 15, 'lutff_6/in_2')

reg n1208 = 0;
// (17, 15, 'sp12_h_r_0')
// (18, 15, 'sp12_h_r_3')
// (19, 15, 'local_g1_4')
// (19, 15, 'lutff_6/in_3')
// (19, 15, 'sp12_h_r_4')
// (20, 15, 'sp12_h_r_7')
// (21, 15, 'sp12_h_r_8')
// (22, 14, 'neigh_op_tnr_2')
// (22, 15, 'neigh_op_rgt_2')
// (22, 15, 'sp12_h_r_11')
// (22, 16, 'neigh_op_bnr_2')
// (23, 14, 'neigh_op_top_2')
// (23, 15, 'lutff_2/out')
// (23, 15, 'sp12_h_r_12')
// (23, 16, 'neigh_op_bot_2')
// (24, 14, 'neigh_op_tnl_2')
// (24, 15, 'neigh_op_lft_2')
// (24, 15, 'sp12_h_r_15')
// (24, 16, 'neigh_op_bnl_2')
// (25, 15, 'sp12_h_r_16')
// (26, 15, 'sp12_h_r_19')
// (27, 15, 'sp12_h_r_20')
// (28, 15, 'sp12_h_r_23')
// (29, 15, 'sp12_h_l_23')

reg n1209 = 0;
// (17, 16, 'local_g0_1')
// (17, 16, 'lutff_2/in_1')
// (17, 16, 'sp4_h_r_9')
// (18, 16, 'sp4_h_r_20')
// (19, 16, 'sp4_h_r_33')
// (20, 13, 'sp4_r_v_b_44')
// (20, 14, 'sp4_r_v_b_33')
// (20, 15, 'sp4_r_v_b_20')
// (20, 16, 'sp4_h_r_44')
// (20, 16, 'sp4_r_v_b_9')
// (21, 11, 'neigh_op_tnr_7')
// (21, 12, 'neigh_op_rgt_7')
// (21, 12, 'sp4_h_r_3')
// (21, 12, 'sp4_v_t_44')
// (21, 13, 'neigh_op_bnr_7')
// (21, 13, 'sp4_v_b_44')
// (21, 14, 'sp4_v_b_33')
// (21, 15, 'sp4_v_b_20')
// (21, 16, 'sp4_h_l_44')
// (21, 16, 'sp4_v_b_9')
// (22, 11, 'neigh_op_top_7')
// (22, 12, 'lutff_7/out')
// (22, 12, 'sp4_h_r_14')
// (22, 13, 'neigh_op_bot_7')
// (23, 11, 'neigh_op_tnl_7')
// (23, 12, 'neigh_op_lft_7')
// (23, 12, 'sp4_h_r_27')
// (23, 13, 'neigh_op_bnl_7')
// (24, 12, 'sp4_h_r_38')
// (25, 12, 'sp4_h_l_38')

reg n1210 = 0;
// (17, 16, 'local_g1_1')
// (17, 16, 'lutff_0/in_0')
// (17, 16, 'sp4_h_r_1')
// (18, 16, 'sp4_h_r_12')
// (19, 16, 'sp4_h_r_25')
// (20, 16, 'sp4_h_r_36')
// (21, 16, 'sp4_h_l_36')
// (21, 16, 'sp4_h_r_1')
// (22, 16, 'sp4_h_r_12')
// (23, 15, 'neigh_op_tnr_2')
// (23, 16, 'neigh_op_rgt_2')
// (23, 16, 'sp4_h_r_25')
// (23, 17, 'neigh_op_bnr_2')
// (24, 15, 'neigh_op_top_2')
// (24, 16, 'lutff_2/out')
// (24, 16, 'sp4_h_r_36')
// (24, 17, 'neigh_op_bot_2')
// (25, 15, 'neigh_op_tnl_2')
// (25, 16, 'neigh_op_lft_2')
// (25, 16, 'sp4_h_l_36')
// (25, 17, 'neigh_op_bnl_2')

reg n1211 = 0;
// (17, 16, 'local_g1_3')
// (17, 16, 'lutff_4/in_0')
// (17, 16, 'sp4_h_r_11')
// (18, 16, 'sp4_h_r_22')
// (19, 15, 'neigh_op_tnr_7')
// (19, 16, 'neigh_op_rgt_7')
// (19, 16, 'sp4_h_r_35')
// (19, 17, 'neigh_op_bnr_7')
// (20, 15, 'neigh_op_top_7')
// (20, 16, 'lutff_7/out')
// (20, 16, 'sp4_h_r_46')
// (20, 17, 'neigh_op_bot_7')
// (21, 15, 'neigh_op_tnl_7')
// (21, 16, 'neigh_op_lft_7')
// (21, 16, 'sp4_h_l_46')
// (21, 17, 'neigh_op_bnl_7')

wire n1212;
// (17, 16, 'lutff_2/lout')
// (17, 16, 'lutff_3/in_2')

wire n1213;
// (17, 16, 'lutff_4/lout')
// (17, 16, 'lutff_5/in_2')

wire n1214;
// (17, 16, 'lutff_5/lout')
// (17, 16, 'lutff_6/in_2')

wire n1215;
// (17, 16, 'neigh_op_tnr_0')
// (17, 17, 'neigh_op_rgt_0')
// (17, 18, 'neigh_op_bnr_0')
// (18, 16, 'neigh_op_top_0')
// (18, 17, 'local_g1_0')
// (18, 17, 'lutff_0/out')
// (18, 17, 'lutff_2/in_1')
// (18, 18, 'neigh_op_bot_0')
// (19, 16, 'neigh_op_tnl_0')
// (19, 17, 'neigh_op_lft_0')
// (19, 18, 'neigh_op_bnl_0')

reg n1216 = 0;
// (17, 16, 'neigh_op_tnr_3')
// (17, 17, 'neigh_op_rgt_3')
// (17, 18, 'neigh_op_bnr_3')
// (18, 16, 'neigh_op_top_3')
// (18, 17, 'local_g1_3')
// (18, 17, 'lutff_1/in_3')
// (18, 17, 'lutff_3/out')
// (18, 18, 'neigh_op_bot_3')
// (19, 16, 'neigh_op_tnl_3')
// (19, 17, 'neigh_op_lft_3')
// (19, 18, 'neigh_op_bnl_3')

wire n1217;
// (17, 16, 'neigh_op_tnr_6')
// (17, 17, 'neigh_op_rgt_6')
// (17, 18, 'neigh_op_bnr_6')
// (18, 11, 'sp12_v_t_23')
// (18, 12, 'sp12_v_b_23')
// (18, 13, 'sp12_v_b_20')
// (18, 14, 'local_g3_3')
// (18, 14, 'lutff_0/in_0')
// (18, 14, 'sp12_v_b_19')
// (18, 15, 'sp12_v_b_16')
// (18, 16, 'neigh_op_top_6')
// (18, 16, 'sp12_v_b_15')
// (18, 17, 'lutff_6/out')
// (18, 17, 'sp12_v_b_12')
// (18, 18, 'neigh_op_bot_6')
// (18, 18, 'sp12_v_b_11')
// (18, 19, 'sp12_v_b_8')
// (18, 20, 'sp12_v_b_7')
// (18, 21, 'sp12_v_b_4')
// (18, 22, 'sp12_v_b_3')
// (18, 23, 'sp12_v_b_0')
// (19, 16, 'neigh_op_tnl_6')
// (19, 17, 'neigh_op_lft_6')
// (19, 18, 'neigh_op_bnl_6')

wire n1218;
// (17, 16, 'neigh_op_tnr_7')
// (17, 17, 'neigh_op_rgt_7')
// (17, 18, 'neigh_op_bnr_7')
// (18, 16, 'neigh_op_top_7')
// (18, 17, 'local_g1_7')
// (18, 17, 'lutff_5/in_3')
// (18, 17, 'lutff_7/out')
// (18, 18, 'neigh_op_bot_7')
// (19, 16, 'neigh_op_tnl_7')
// (19, 17, 'neigh_op_lft_7')
// (19, 18, 'neigh_op_bnl_7')

reg n1219 = 0;
// (17, 17, 'local_g0_6')
// (17, 17, 'lutff_5/in_1')
// (17, 17, 'sp4_h_r_6')
// (18, 17, 'sp4_h_r_19')
// (19, 17, 'sp4_h_r_30')
// (20, 17, 'sp4_h_r_43')
// (21, 17, 'sp4_h_l_43')
// (21, 17, 'sp4_h_r_6')
// (22, 17, 'sp4_h_r_19')
// (23, 17, 'neigh_op_tnr_2')
// (23, 17, 'sp4_h_r_30')
// (23, 18, 'neigh_op_rgt_2')
// (23, 19, 'neigh_op_bnr_2')
// (24, 17, 'neigh_op_top_2')
// (24, 17, 'sp4_h_r_43')
// (24, 18, 'lutff_2/out')
// (24, 18, 'sp4_r_v_b_37')
// (24, 19, 'neigh_op_bot_2')
// (24, 19, 'sp4_r_v_b_24')
// (24, 20, 'sp4_r_v_b_13')
// (24, 21, 'sp4_r_v_b_0')
// (25, 17, 'neigh_op_tnl_2')
// (25, 17, 'sp4_h_l_43')
// (25, 17, 'sp4_v_t_37')
// (25, 18, 'neigh_op_lft_2')
// (25, 18, 'sp4_v_b_37')
// (25, 19, 'neigh_op_bnl_2')
// (25, 19, 'sp4_v_b_24')
// (25, 20, 'sp4_v_b_13')
// (25, 21, 'sp4_v_b_0')

wire n1220;
// (17, 17, 'lutff_1/lout')
// (17, 17, 'lutff_2/in_2')

wire n1221;
// (17, 17, 'lutff_5/lout')
// (17, 17, 'lutff_6/in_2')

wire n1222;
// (17, 17, 'neigh_op_tnr_0')
// (17, 18, 'neigh_op_rgt_0')
// (17, 19, 'neigh_op_bnr_0')
// (18, 17, 'neigh_op_top_0')
// (18, 18, 'local_g3_0')
// (18, 18, 'lutff_0/out')
// (18, 18, 'lutff_2/in_1')
// (18, 19, 'neigh_op_bot_0')
// (19, 17, 'neigh_op_tnl_0')
// (19, 18, 'neigh_op_lft_0')
// (19, 19, 'neigh_op_bnl_0')

wire n1223;
// (17, 17, 'neigh_op_tnr_2')
// (17, 18, 'neigh_op_rgt_2')
// (17, 19, 'neigh_op_bnr_2')
// (18, 17, 'neigh_op_top_2')
// (18, 18, 'lutff_2/out')
// (18, 19, 'neigh_op_bot_2')
// (19, 17, 'local_g3_2')
// (19, 17, 'lutff_6/in_3')
// (19, 17, 'neigh_op_tnl_2')
// (19, 18, 'neigh_op_lft_2')
// (19, 19, 'neigh_op_bnl_2')

reg n1224 = 0;
// (17, 17, 'neigh_op_tnr_3')
// (17, 18, 'neigh_op_rgt_3')
// (17, 19, 'neigh_op_bnr_3')
// (18, 17, 'neigh_op_top_3')
// (18, 18, 'local_g3_3')
// (18, 18, 'lutff_1/in_3')
// (18, 18, 'lutff_3/out')
// (18, 19, 'neigh_op_bot_3')
// (19, 17, 'neigh_op_tnl_3')
// (19, 18, 'neigh_op_lft_3')
// (19, 19, 'neigh_op_bnl_3')

wire n1225;
// (17, 17, 'neigh_op_tnr_4')
// (17, 18, 'neigh_op_rgt_4')
// (17, 19, 'neigh_op_bnr_4')
// (18, 17, 'neigh_op_top_4')
// (18, 18, 'local_g1_4')
// (18, 18, 'lutff_4/out')
// (18, 18, 'lutff_6/in_3')
// (18, 19, 'neigh_op_bot_4')
// (19, 17, 'neigh_op_tnl_4')
// (19, 18, 'neigh_op_lft_4')
// (19, 19, 'neigh_op_bnl_4')

reg n1226 = 0;
// (17, 17, 'sp12_h_r_1')
// (18, 17, 'sp12_h_r_2')
// (19, 17, 'sp12_h_r_5')
// (20, 17, 'local_g1_6')
// (20, 17, 'lutff_6/in_1')
// (20, 17, 'sp12_h_r_6')
// (21, 17, 'sp12_h_r_9')
// (22, 17, 'sp12_h_r_10')
// (23, 16, 'neigh_op_tnr_3')
// (23, 17, 'neigh_op_rgt_3')
// (23, 17, 'sp12_h_r_13')
// (23, 18, 'neigh_op_bnr_3')
// (24, 16, 'neigh_op_top_3')
// (24, 17, 'lutff_3/out')
// (24, 17, 'sp12_h_r_14')
// (24, 18, 'neigh_op_bot_3')
// (25, 16, 'neigh_op_tnl_3')
// (25, 17, 'neigh_op_lft_3')
// (25, 17, 'sp12_h_r_17')
// (25, 18, 'neigh_op_bnl_3')
// (26, 17, 'sp12_h_r_18')
// (27, 17, 'sp12_h_r_21')
// (28, 17, 'sp12_h_r_22')
// (29, 17, 'sp12_h_l_22')

reg n1227 = 0;
// (17, 17, 'sp4_h_r_8')
// (18, 17, 'local_g1_5')
// (18, 17, 'lutff_1/in_1')
// (18, 17, 'sp4_h_r_21')
// (19, 17, 'sp4_h_r_32')
// (20, 17, 'sp4_h_r_45')
// (20, 18, 'sp4_r_v_b_45')
// (20, 19, 'sp4_r_v_b_32')
// (20, 20, 'sp4_r_v_b_21')
// (20, 21, 'sp4_r_v_b_8')
// (21, 17, 'sp4_h_l_45')
// (21, 17, 'sp4_v_t_45')
// (21, 18, 'sp4_v_b_45')
// (21, 19, 'sp4_v_b_32')
// (21, 20, 'neigh_op_tnr_7')
// (21, 20, 'sp4_v_b_21')
// (21, 21, 'neigh_op_rgt_7')
// (21, 21, 'sp4_h_r_3')
// (21, 21, 'sp4_v_b_8')
// (21, 22, 'neigh_op_bnr_7')
// (22, 20, 'neigh_op_top_7')
// (22, 21, 'lutff_7/out')
// (22, 21, 'sp4_h_r_14')
// (22, 22, 'neigh_op_bot_7')
// (23, 20, 'neigh_op_tnl_7')
// (23, 21, 'neigh_op_lft_7')
// (23, 21, 'sp4_h_r_27')
// (23, 22, 'neigh_op_bnl_7')
// (24, 21, 'sp4_h_r_38')
// (25, 21, 'sp4_h_l_38')

reg n1228 = 0;
// (17, 17, 'sp4_r_v_b_36')
// (17, 18, 'sp4_r_v_b_25')
// (17, 19, 'sp4_r_v_b_12')
// (17, 20, 'sp4_r_v_b_1')
// (18, 16, 'sp4_v_t_36')
// (18, 17, 'sp4_v_b_36')
// (18, 18, 'sp4_v_b_25')
// (18, 19, 'local_g0_4')
// (18, 19, 'lutff_5/in_1')
// (18, 19, 'sp4_v_b_12')
// (18, 20, 'sp4_h_r_1')
// (18, 20, 'sp4_v_b_1')
// (19, 20, 'sp4_h_r_12')
// (20, 20, 'sp4_h_r_25')
// (21, 20, 'sp4_h_r_36')
// (22, 19, 'neigh_op_tnr_0')
// (22, 20, 'neigh_op_rgt_0')
// (22, 20, 'sp4_h_l_36')
// (22, 20, 'sp4_h_r_5')
// (22, 21, 'neigh_op_bnr_0')
// (23, 19, 'neigh_op_top_0')
// (23, 20, 'lutff_0/out')
// (23, 20, 'sp4_h_r_16')
// (23, 21, 'neigh_op_bot_0')
// (24, 19, 'neigh_op_tnl_0')
// (24, 20, 'neigh_op_lft_0')
// (24, 20, 'sp4_h_r_29')
// (24, 21, 'neigh_op_bnl_0')
// (25, 20, 'sp4_h_r_40')
// (26, 20, 'sp4_h_l_40')

reg n1229 = 0;
// (17, 17, 'sp4_r_v_b_37')
// (17, 18, 'sp4_r_v_b_24')
// (17, 19, 'sp4_r_v_b_13')
// (17, 20, 'sp4_r_v_b_0')
// (18, 16, 'sp4_v_t_37')
// (18, 17, 'sp4_v_b_37')
// (18, 18, 'sp4_v_b_24')
// (18, 19, 'local_g0_5')
// (18, 19, 'lutff_6/in_1')
// (18, 19, 'sp4_v_b_13')
// (18, 20, 'sp4_h_r_7')
// (18, 20, 'sp4_v_b_0')
// (19, 20, 'sp4_h_r_18')
// (20, 20, 'sp4_h_r_31')
// (21, 20, 'sp4_h_r_42')
// (22, 19, 'neigh_op_tnr_1')
// (22, 20, 'neigh_op_rgt_1')
// (22, 20, 'sp4_h_l_42')
// (22, 20, 'sp4_h_r_7')
// (22, 21, 'neigh_op_bnr_1')
// (23, 19, 'neigh_op_top_1')
// (23, 20, 'lutff_1/out')
// (23, 20, 'sp4_h_r_18')
// (23, 21, 'neigh_op_bot_1')
// (24, 19, 'neigh_op_tnl_1')
// (24, 20, 'neigh_op_lft_1')
// (24, 20, 'sp4_h_r_31')
// (24, 21, 'neigh_op_bnl_1')
// (25, 20, 'sp4_h_r_42')
// (26, 20, 'sp4_h_l_42')

wire n1230;
// (17, 17, 'sp4_r_v_b_44')
// (17, 18, 'neigh_op_tnr_2')
// (17, 18, 'sp4_r_v_b_33')
// (17, 19, 'neigh_op_rgt_2')
// (17, 19, 'sp4_r_v_b_20')
// (17, 20, 'neigh_op_bnr_2')
// (17, 20, 'sp4_r_v_b_9')
// (18, 16, 'sp4_v_t_44')
// (18, 17, 'local_g3_4')
// (18, 17, 'lutff_6/in_1')
// (18, 17, 'sp4_v_b_44')
// (18, 18, 'neigh_op_top_2')
// (18, 18, 'sp4_v_b_33')
// (18, 19, 'lutff_2/out')
// (18, 19, 'sp4_v_b_20')
// (18, 20, 'neigh_op_bot_2')
// (18, 20, 'sp4_v_b_9')
// (19, 18, 'neigh_op_tnl_2')
// (19, 19, 'neigh_op_lft_2')
// (19, 20, 'neigh_op_bnl_2')

wire n1231;
// (17, 18, 'lutff_7/cout')
// (17, 19, 'carry_in')
// (17, 19, 'carry_in_mux')

wire n1232;
// (17, 18, 'neigh_op_tnr_0')
// (17, 19, 'neigh_op_rgt_0')
// (17, 20, 'neigh_op_bnr_0')
// (18, 18, 'local_g0_0')
// (18, 18, 'lutff_7/in_1')
// (18, 18, 'neigh_op_top_0')
// (18, 19, 'lutff_0/out')
// (18, 20, 'neigh_op_bot_0')
// (19, 18, 'neigh_op_tnl_0')
// (19, 19, 'neigh_op_lft_0')
// (19, 20, 'neigh_op_bnl_0')

reg n1233 = 0;
// (17, 18, 'neigh_op_tnr_1')
// (17, 19, 'neigh_op_rgt_1')
// (17, 20, 'neigh_op_bnr_1')
// (18, 18, 'neigh_op_top_1')
// (18, 19, 'local_g2_1')
// (18, 19, 'lutff_0/in_3')
// (18, 19, 'lutff_1/out')
// (18, 20, 'neigh_op_bot_1')
// (19, 18, 'neigh_op_tnl_1')
// (19, 19, 'neigh_op_lft_1')
// (19, 20, 'neigh_op_bnl_1')

wire n1234;
// (17, 18, 'neigh_op_tnr_3')
// (17, 19, 'neigh_op_rgt_3')
// (17, 20, 'neigh_op_bnr_3')
// (18, 17, 'sp4_r_v_b_47')
// (18, 18, 'neigh_op_top_3')
// (18, 18, 'sp4_r_v_b_34')
// (18, 19, 'lutff_3/out')
// (18, 19, 'sp4_r_v_b_23')
// (18, 20, 'neigh_op_bot_3')
// (18, 20, 'sp4_r_v_b_10')
// (19, 16, 'sp4_v_t_47')
// (19, 17, 'sp4_v_b_47')
// (19, 18, 'neigh_op_tnl_3')
// (19, 18, 'sp4_v_b_34')
// (19, 19, 'neigh_op_lft_3')
// (19, 19, 'sp4_v_b_23')
// (19, 20, 'neigh_op_bnl_3')
// (19, 20, 'sp4_h_r_4')
// (19, 20, 'sp4_v_b_10')
// (20, 20, 'sp4_h_r_17')
// (21, 20, 'sp4_h_r_28')
// (22, 20, 'local_g3_1')
// (22, 20, 'lutff_4/in_0')
// (22, 20, 'sp4_h_r_41')
// (23, 20, 'sp4_h_l_41')

wire n1235;
// (17, 18, 'neigh_op_tnr_4')
// (17, 19, 'neigh_op_rgt_4')
// (17, 20, 'neigh_op_bnr_4')
// (18, 18, 'local_g0_4')
// (18, 18, 'lutff_7/in_3')
// (18, 18, 'neigh_op_top_4')
// (18, 19, 'lutff_4/out')
// (18, 20, 'neigh_op_bot_4')
// (19, 18, 'neigh_op_tnl_4')
// (19, 19, 'neigh_op_lft_4')
// (19, 20, 'neigh_op_bnl_4')

wire n1236;
// (17, 18, 'neigh_op_tnr_5')
// (17, 19, 'neigh_op_rgt_5')
// (17, 20, 'neigh_op_bnr_5')
// (18, 12, 'sp12_v_t_22')
// (18, 13, 'sp12_v_b_22')
// (18, 14, 'local_g3_5')
// (18, 14, 'lutff_4/in_0')
// (18, 14, 'sp12_v_b_21')
// (18, 15, 'sp12_v_b_18')
// (18, 16, 'sp12_v_b_17')
// (18, 17, 'sp12_v_b_14')
// (18, 18, 'neigh_op_top_5')
// (18, 18, 'sp12_v_b_13')
// (18, 19, 'lutff_5/out')
// (18, 19, 'sp12_v_b_10')
// (18, 20, 'neigh_op_bot_5')
// (18, 20, 'sp12_v_b_9')
// (18, 21, 'sp12_v_b_6')
// (18, 22, 'sp12_v_b_5')
// (18, 23, 'sp12_v_b_2')
// (18, 24, 'sp12_v_b_1')
// (19, 18, 'neigh_op_tnl_5')
// (19, 19, 'neigh_op_lft_5')
// (19, 20, 'neigh_op_bnl_5')

wire n1237;
// (17, 18, 'neigh_op_tnr_6')
// (17, 19, 'neigh_op_rgt_6')
// (17, 20, 'neigh_op_bnr_6')
// (18, 15, 'sp4_r_v_b_45')
// (18, 16, 'sp4_r_v_b_32')
// (18, 17, 'sp4_r_v_b_21')
// (18, 18, 'neigh_op_top_6')
// (18, 18, 'sp4_r_v_b_8')
// (18, 19, 'lutff_6/out')
// (18, 19, 'sp4_r_v_b_45')
// (18, 20, 'neigh_op_bot_6')
// (18, 20, 'sp4_r_v_b_32')
// (18, 21, 'sp4_r_v_b_21')
// (18, 22, 'sp4_r_v_b_8')
// (19, 14, 'sp4_h_r_1')
// (19, 14, 'sp4_v_t_45')
// (19, 15, 'sp4_v_b_45')
// (19, 16, 'sp4_v_b_32')
// (19, 17, 'sp4_v_b_21')
// (19, 18, 'neigh_op_tnl_6')
// (19, 18, 'sp4_v_b_8')
// (19, 18, 'sp4_v_t_45')
// (19, 19, 'neigh_op_lft_6')
// (19, 19, 'sp4_v_b_45')
// (19, 20, 'neigh_op_bnl_6')
// (19, 20, 'sp4_v_b_32')
// (19, 21, 'sp4_v_b_21')
// (19, 22, 'sp4_v_b_8')
// (20, 14, 'local_g0_4')
// (20, 14, 'lutff_3/in_3')
// (20, 14, 'sp4_h_r_12')
// (21, 14, 'sp4_h_r_25')
// (22, 14, 'sp4_h_r_36')
// (23, 14, 'sp4_h_l_36')

reg n1238 = 0;
// (17, 18, 'sp4_h_r_5')
// (18, 18, 'sp4_h_r_16')
// (19, 17, 'neigh_op_tnr_4')
// (19, 18, 'neigh_op_rgt_4')
// (19, 18, 'sp4_h_r_29')
// (19, 19, 'neigh_op_bnr_4')
// (20, 17, 'neigh_op_top_4')
// (20, 18, 'lutff_4/out')
// (20, 18, 'sp4_h_r_40')
// (20, 19, 'neigh_op_bot_4')
// (20, 19, 'sp4_r_v_b_40')
// (20, 20, 'sp4_r_v_b_29')
// (20, 21, 'sp4_r_v_b_16')
// (20, 22, 'sp4_r_v_b_5')
// (21, 17, 'neigh_op_tnl_4')
// (21, 18, 'neigh_op_lft_4')
// (21, 18, 'sp4_h_l_40')
// (21, 18, 'sp4_v_t_40')
// (21, 19, 'neigh_op_bnl_4')
// (21, 19, 'sp4_v_b_40')
// (21, 20, 'sp4_v_b_29')
// (21, 21, 'sp4_v_b_16')
// (21, 22, 'local_g0_5')
// (21, 22, 'lutff_2/in_3')
// (21, 22, 'sp4_v_b_5')

wire n1239;
// (17, 18, 'sp4_r_v_b_38')
// (17, 19, 'neigh_op_tnr_7')
// (17, 19, 'sp4_r_v_b_27')
// (17, 20, 'neigh_op_rgt_7')
// (17, 20, 'sp4_r_v_b_14')
// (17, 21, 'neigh_op_bnr_7')
// (17, 21, 'sp4_r_v_b_3')
// (18, 17, 'sp4_v_t_38')
// (18, 18, 'local_g3_6')
// (18, 18, 'lutff_2/in_3')
// (18, 18, 'sp4_v_b_38')
// (18, 19, 'neigh_op_top_7')
// (18, 19, 'sp4_v_b_27')
// (18, 20, 'lutff_7/out')
// (18, 20, 'sp4_v_b_14')
// (18, 21, 'neigh_op_bot_7')
// (18, 21, 'sp4_v_b_3')
// (19, 19, 'neigh_op_tnl_7')
// (19, 20, 'neigh_op_lft_7')
// (19, 21, 'neigh_op_bnl_7')

reg n1240 = 0;
// (17, 18, 'sp4_r_v_b_41')
// (17, 19, 'sp4_r_v_b_28')
// (17, 20, 'sp4_r_v_b_17')
// (17, 21, 'local_g1_4')
// (17, 21, 'lutff_6/in_1')
// (17, 21, 'sp4_r_v_b_4')
// (18, 17, 'sp4_h_r_10')
// (18, 17, 'sp4_v_t_41')
// (18, 18, 'sp4_v_b_41')
// (18, 19, 'sp4_v_b_28')
// (18, 20, 'sp4_v_b_17')
// (18, 21, 'sp4_v_b_4')
// (19, 17, 'sp4_h_r_23')
// (20, 17, 'sp4_h_r_34')
// (21, 17, 'sp4_h_r_47')
// (22, 17, 'sp4_h_l_47')
// (22, 17, 'sp4_h_r_2')
// (23, 16, 'neigh_op_tnr_5')
// (23, 17, 'neigh_op_rgt_5')
// (23, 17, 'sp4_h_r_15')
// (23, 18, 'neigh_op_bnr_5')
// (24, 16, 'neigh_op_top_5')
// (24, 17, 'lutff_5/out')
// (24, 17, 'sp4_h_r_26')
// (24, 18, 'neigh_op_bot_5')
// (25, 16, 'neigh_op_tnl_5')
// (25, 17, 'neigh_op_lft_5')
// (25, 17, 'sp4_h_r_39')
// (25, 18, 'neigh_op_bnl_5')
// (26, 17, 'sp4_h_l_39')

wire n1241;
// (17, 18, 'sp4_r_v_b_43')
// (17, 19, 'sp4_r_v_b_30')
// (17, 20, 'sp4_r_v_b_19')
// (17, 21, 'sp4_r_v_b_6')
// (17, 22, 'sp4_r_v_b_38')
// (17, 23, 'neigh_op_tnr_7')
// (17, 23, 'sp4_r_v_b_27')
// (17, 24, 'neigh_op_rgt_7')
// (17, 24, 'sp4_r_v_b_14')
// (17, 25, 'neigh_op_bnr_7')
// (17, 25, 'sp4_r_v_b_3')
// (18, 17, 'local_g1_6')
// (18, 17, 'lutff_2/in_3')
// (18, 17, 'sp4_h_r_6')
// (18, 17, 'sp4_v_t_43')
// (18, 18, 'sp4_v_b_43')
// (18, 19, 'sp4_v_b_30')
// (18, 20, 'sp4_v_b_19')
// (18, 21, 'sp4_v_b_6')
// (18, 21, 'sp4_v_t_38')
// (18, 22, 'sp4_v_b_38')
// (18, 23, 'neigh_op_top_7')
// (18, 23, 'sp4_v_b_27')
// (18, 24, 'lutff_7/out')
// (18, 24, 'sp4_v_b_14')
// (18, 25, 'neigh_op_bot_7')
// (18, 25, 'sp4_v_b_3')
// (19, 17, 'sp4_h_r_19')
// (19, 23, 'neigh_op_tnl_7')
// (19, 24, 'neigh_op_lft_7')
// (19, 25, 'neigh_op_bnl_7')
// (20, 17, 'sp4_h_r_30')
// (21, 17, 'sp4_h_r_43')
// (22, 17, 'sp4_h_l_43')

wire n1242;
// (17, 18, 'sp4_r_v_b_45')
// (17, 19, 'sp4_r_v_b_32')
// (17, 20, 'sp4_r_v_b_21')
// (17, 21, 'sp4_r_v_b_8')
// (18, 17, 'sp12_v_t_23')
// (18, 17, 'sp4_v_t_45')
// (18, 18, 'sp12_v_b_23')
// (18, 18, 'sp4_v_b_45')
// (18, 19, 'sp12_v_b_20')
// (18, 19, 'sp4_v_b_32')
// (18, 20, 'sp12_v_b_19')
// (18, 20, 'sp4_v_b_21')
// (18, 21, 'sp12_v_b_16')
// (18, 21, 'sp4_h_r_8')
// (18, 21, 'sp4_v_b_8')
// (18, 22, 'sp12_v_b_15')
// (18, 23, 'sp12_v_b_12')
// (18, 24, 'sp12_v_b_11')
// (18, 25, 'sp12_v_b_8')
// (18, 26, 'sp12_v_b_7')
// (18, 27, 'sp12_v_b_4')
// (18, 28, 'sp12_v_b_3')
// (18, 29, 'sp12_h_r_0')
// (18, 29, 'sp12_v_b_0')
// (19, 21, 'local_g1_5')
// (19, 21, 'lutff_4/in_2')
// (19, 21, 'sp4_h_r_21')
// (19, 29, 'sp12_h_r_3')
// (20, 21, 'sp4_h_r_32')
// (20, 29, 'sp12_h_r_4')
// (21, 21, 'sp4_h_r_45')
// (21, 29, 'sp12_h_r_7')
// (22, 21, 'sp4_h_l_45')
// (22, 29, 'sp12_h_r_8')
// (23, 29, 'sp12_h_r_11')
// (24, 29, 'sp12_h_r_12')
// (25, 29, 'sp12_h_r_15')
// (26, 29, 'sp12_h_r_16')
// (27, 29, 'sp12_h_r_19')
// (28, 29, 'sp12_h_r_20')
// (29, 29, 'sp12_h_r_23')
// (29, 32, 'neigh_op_tnr_0')
// (29, 32, 'neigh_op_tnr_4')
// (30, 29, 'sp12_h_l_23')
// (30, 29, 'sp12_v_t_23')
// (30, 30, 'sp12_v_b_23')
// (30, 31, 'sp12_v_b_20')
// (30, 32, 'neigh_op_top_0')
// (30, 32, 'neigh_op_top_4')
// (30, 32, 'sp12_v_b_19')
// (30, 33, 'io_0/D_IN_0')
// (30, 33, 'span12_vert_16')
// (31, 32, 'neigh_op_tnl_0')
// (31, 32, 'neigh_op_tnl_4')

reg n1243 = 0;
// (17, 18, 'sp4_r_v_b_46')
// (17, 19, 'sp4_r_v_b_35')
// (17, 20, 'sp4_r_v_b_22')
// (17, 21, 'local_g2_3')
// (17, 21, 'lutff_6/in_3')
// (17, 21, 'sp4_r_v_b_11')
// (18, 17, 'sp4_h_r_5')
// (18, 17, 'sp4_v_t_46')
// (18, 18, 'sp4_v_b_46')
// (18, 19, 'sp4_v_b_35')
// (18, 20, 'sp4_v_b_22')
// (18, 21, 'sp4_v_b_11')
// (19, 17, 'sp4_h_r_16')
// (20, 17, 'sp4_h_r_29')
// (21, 14, 'sp4_r_v_b_40')
// (21, 15, 'sp4_r_v_b_29')
// (21, 16, 'sp4_r_v_b_16')
// (21, 17, 'sp4_h_r_40')
// (21, 17, 'sp4_r_v_b_5')
// (22, 12, 'neigh_op_tnr_3')
// (22, 13, 'neigh_op_rgt_3')
// (22, 13, 'sp4_h_r_11')
// (22, 13, 'sp4_v_t_40')
// (22, 14, 'neigh_op_bnr_3')
// (22, 14, 'sp4_v_b_40')
// (22, 15, 'sp4_v_b_29')
// (22, 16, 'sp4_v_b_16')
// (22, 17, 'sp4_h_l_40')
// (22, 17, 'sp4_v_b_5')
// (23, 12, 'neigh_op_top_3')
// (23, 13, 'lutff_3/out')
// (23, 13, 'sp4_h_r_22')
// (23, 14, 'neigh_op_bot_3')
// (24, 12, 'neigh_op_tnl_3')
// (24, 13, 'neigh_op_lft_3')
// (24, 13, 'sp4_h_r_35')
// (24, 14, 'neigh_op_bnl_3')
// (25, 13, 'sp4_h_r_46')
// (26, 13, 'sp4_h_l_46')

wire n1244;
// (17, 19, 'lutff_7/cout')
// (17, 20, 'carry_in')
// (17, 20, 'carry_in_mux')

wire n1245;
// (17, 19, 'neigh_op_tnr_2')
// (17, 20, 'neigh_op_rgt_2')
// (17, 21, 'neigh_op_bnr_2')
// (18, 19, 'neigh_op_top_2')
// (18, 20, 'lutff_2/out')
// (18, 20, 'sp4_h_r_4')
// (18, 21, 'neigh_op_bot_2')
// (19, 19, 'neigh_op_tnl_2')
// (19, 20, 'neigh_op_lft_2')
// (19, 20, 'sp4_h_r_17')
// (19, 21, 'neigh_op_bnl_2')
// (20, 20, 'sp4_h_r_28')
// (21, 17, 'sp4_r_v_b_47')
// (21, 18, 'sp4_r_v_b_34')
// (21, 19, 'sp4_r_v_b_23')
// (21, 20, 'sp4_h_r_41')
// (21, 20, 'sp4_r_v_b_10')
// (22, 16, 'sp4_v_t_47')
// (22, 17, 'sp4_v_b_47')
// (22, 18, 'local_g3_2')
// (22, 18, 'lutff_6/in_3')
// (22, 18, 'sp4_v_b_34')
// (22, 19, 'sp4_v_b_23')
// (22, 20, 'sp4_h_l_41')
// (22, 20, 'sp4_v_b_10')

wire n1246;
// (17, 19, 'neigh_op_tnr_4')
// (17, 20, 'neigh_op_rgt_4')
// (17, 21, 'neigh_op_bnr_4')
// (18, 19, 'neigh_op_top_4')
// (18, 20, 'local_g1_4')
// (18, 20, 'lutff_2/in_3')
// (18, 20, 'lutff_4/out')
// (18, 21, 'neigh_op_bot_4')
// (19, 19, 'neigh_op_tnl_4')
// (19, 20, 'neigh_op_lft_4')
// (19, 21, 'neigh_op_bnl_4')

wire n1247;
// (17, 19, 'neigh_op_tnr_5')
// (17, 20, 'neigh_op_rgt_5')
// (17, 21, 'neigh_op_bnr_5')
// (18, 19, 'neigh_op_top_5')
// (18, 20, 'local_g2_5')
// (18, 20, 'lutff_2/in_1')
// (18, 20, 'lutff_5/out')
// (18, 21, 'neigh_op_bot_5')
// (19, 19, 'neigh_op_tnl_5')
// (19, 20, 'neigh_op_lft_5')
// (19, 21, 'neigh_op_bnl_5')

reg n1248 = 0;
// (17, 19, 'neigh_op_tnr_6')
// (17, 20, 'neigh_op_rgt_6')
// (17, 21, 'neigh_op_bnr_6')
// (18, 19, 'neigh_op_top_6')
// (18, 20, 'local_g3_6')
// (18, 20, 'lutff_0/in_3')
// (18, 20, 'lutff_6/out')
// (18, 21, 'neigh_op_bot_6')
// (19, 19, 'neigh_op_tnl_6')
// (19, 20, 'neigh_op_lft_6')
// (19, 21, 'neigh_op_bnl_6')

reg n1249 = 0;
// (17, 19, 'sp4_h_r_3')
// (18, 19, 'local_g0_6')
// (18, 19, 'lutff_3/in_3')
// (18, 19, 'sp4_h_r_14')
// (19, 18, 'neigh_op_tnr_3')
// (19, 19, 'neigh_op_rgt_3')
// (19, 19, 'sp4_h_r_27')
// (19, 20, 'neigh_op_bnr_3')
// (20, 18, 'neigh_op_top_3')
// (20, 19, 'lutff_3/out')
// (20, 19, 'sp4_h_r_38')
// (20, 20, 'neigh_op_bot_3')
// (21, 18, 'neigh_op_tnl_3')
// (21, 19, 'neigh_op_lft_3')
// (21, 19, 'sp4_h_l_38')
// (21, 20, 'neigh_op_bnl_3')

reg n1250 = 0;
// (17, 19, 'sp4_r_v_b_36')
// (17, 20, 'sp4_r_v_b_25')
// (17, 21, 'sp4_r_v_b_12')
// (17, 22, 'sp4_r_v_b_1')
// (18, 18, 'sp4_h_r_7')
// (18, 18, 'sp4_v_t_36')
// (18, 19, 'sp4_v_b_36')
// (18, 20, 'local_g2_1')
// (18, 20, 'lutff_4/in_3')
// (18, 20, 'sp4_v_b_25')
// (18, 21, 'sp4_v_b_12')
// (18, 22, 'sp4_v_b_1')
// (19, 18, 'sp4_h_r_18')
// (20, 18, 'sp4_h_r_31')
// (21, 18, 'sp4_h_r_42')
// (22, 17, 'neigh_op_tnr_3')
// (22, 18, 'neigh_op_rgt_3')
// (22, 18, 'sp4_h_l_42')
// (22, 18, 'sp4_h_r_11')
// (22, 19, 'neigh_op_bnr_3')
// (23, 17, 'neigh_op_top_3')
// (23, 18, 'lutff_3/out')
// (23, 18, 'sp4_h_r_22')
// (23, 19, 'neigh_op_bot_3')
// (24, 17, 'neigh_op_tnl_3')
// (24, 18, 'neigh_op_lft_3')
// (24, 18, 'sp4_h_r_35')
// (24, 19, 'neigh_op_bnl_3')
// (25, 18, 'sp4_h_r_46')
// (26, 18, 'sp4_h_l_46')

wire n1251;
// (17, 20, 'lutff_7/cout')
// (17, 21, 'carry_in')
// (17, 21, 'carry_in_mux')
// (17, 21, 'lutff_0/in_3')

reg io_33_3_1 = 0;
// (17, 20, 'neigh_op_tnr_2')
// (17, 21, 'neigh_op_rgt_2')
// (17, 22, 'neigh_op_bnr_2')
// (18, 7, 'sp12_h_r_0')
// (18, 7, 'sp12_v_t_23')
// (18, 8, 'sp12_v_b_23')
// (18, 9, 'sp12_v_b_20')
// (18, 10, 'sp12_v_b_19')
// (18, 11, 'sp12_v_b_16')
// (18, 12, 'sp12_v_b_15')
// (18, 13, 'sp12_v_b_12')
// (18, 14, 'sp12_v_b_11')
// (18, 15, 'sp12_v_b_8')
// (18, 16, 'sp12_v_b_7')
// (18, 17, 'sp12_v_b_4')
// (18, 18, 'sp12_v_b_3')
// (18, 19, 'sp12_v_b_0')
// (18, 19, 'sp12_v_t_23')
// (18, 20, 'neigh_op_top_2')
// (18, 20, 'sp12_v_b_23')
// (18, 21, 'lutff_2/out')
// (18, 21, 'sp12_v_b_20')
// (18, 22, 'neigh_op_bot_2')
// (18, 22, 'sp12_v_b_19')
// (18, 23, 'sp12_v_b_16')
// (18, 24, 'sp12_v_b_15')
// (18, 25, 'sp12_v_b_12')
// (18, 26, 'sp12_v_b_11')
// (18, 27, 'sp12_v_b_8')
// (18, 28, 'sp12_v_b_7')
// (18, 29, 'sp12_v_b_4')
// (18, 30, 'sp12_v_b_3')
// (18, 31, 'sp12_v_b_0')
// (19, 7, 'sp12_h_r_3')
// (19, 20, 'neigh_op_tnl_2')
// (19, 21, 'neigh_op_lft_2')
// (19, 22, 'neigh_op_bnl_2')
// (20, 7, 'sp12_h_r_4')
// (21, 7, 'sp12_h_r_7')
// (22, 7, 'sp12_h_r_8')
// (23, 7, 'sp12_h_r_11')
// (24, 7, 'sp12_h_r_12')
// (25, 7, 'sp12_h_r_15')
// (25, 7, 'sp4_h_r_9')
// (26, 7, 'sp12_h_r_16')
// (26, 7, 'sp4_h_r_20')
// (27, 7, 'sp12_h_r_19')
// (27, 7, 'sp4_h_r_33')
// (28, 4, 'sp4_r_v_b_38')
// (28, 5, 'sp4_r_v_b_27')
// (28, 6, 'sp4_r_v_b_14')
// (28, 7, 'sp12_h_r_20')
// (28, 7, 'sp4_h_r_44')
// (28, 7, 'sp4_r_v_b_3')
// (29, 3, 'sp4_h_r_8')
// (29, 3, 'sp4_v_t_38')
// (29, 4, 'sp4_v_b_38')
// (29, 5, 'sp4_v_b_27')
// (29, 6, 'sp4_v_b_14')
// (29, 7, 'sp12_h_r_23')
// (29, 7, 'sp4_h_l_44')
// (29, 7, 'sp4_v_b_3')
// (30, 3, 'sp4_h_r_21')
// (30, 7, 'sp12_h_l_23')
// (31, 3, 'sp4_h_r_32')
// (32, 3, 'sp4_h_r_45')
// (33, 3, 'io_1/D_OUT_0')
// (33, 3, 'io_1/PAD')
// (33, 3, 'local_g0_5')
// (33, 3, 'span4_horz_45')

reg io_20_33_1 = 0;
// (17, 20, 'neigh_op_tnr_3')
// (17, 21, 'neigh_op_rgt_3')
// (17, 21, 'sp4_h_r_11')
// (17, 22, 'neigh_op_bnr_3')
// (17, 33, 'span4_horz_r_1')
// (18, 20, 'neigh_op_top_3')
// (18, 21, 'lutff_3/out')
// (18, 21, 'sp4_h_r_22')
// (18, 22, 'neigh_op_bot_3')
// (18, 33, 'span4_horz_r_5')
// (19, 20, 'neigh_op_tnl_3')
// (19, 21, 'neigh_op_lft_3')
// (19, 21, 'sp4_h_r_35')
// (19, 22, 'neigh_op_bnl_3')
// (19, 33, 'span4_horz_r_9')
// (20, 21, 'sp4_h_r_46')
// (20, 22, 'sp4_r_v_b_41')
// (20, 23, 'sp4_r_v_b_28')
// (20, 24, 'sp4_r_v_b_17')
// (20, 25, 'sp4_r_v_b_4')
// (20, 26, 'sp4_r_v_b_41')
// (20, 27, 'sp4_r_v_b_28')
// (20, 28, 'sp4_r_v_b_17')
// (20, 29, 'sp4_r_v_b_4')
// (20, 30, 'sp4_r_v_b_42')
// (20, 31, 'sp4_r_v_b_31')
// (20, 32, 'sp4_r_v_b_18')
// (20, 33, 'io_1/D_OUT_0')
// (20, 33, 'io_1/PAD')
// (20, 33, 'local_g0_5')
// (20, 33, 'span4_horz_r_13')
// (21, 21, 'sp4_h_l_46')
// (21, 21, 'sp4_v_t_41')
// (21, 22, 'sp4_v_b_41')
// (21, 23, 'sp4_v_b_28')
// (21, 24, 'sp4_v_b_17')
// (21, 25, 'sp4_v_b_4')
// (21, 25, 'sp4_v_t_41')
// (21, 26, 'sp4_v_b_41')
// (21, 27, 'sp4_v_b_28')
// (21, 28, 'sp4_v_b_17')
// (21, 29, 'sp4_v_b_4')
// (21, 29, 'sp4_v_t_42')
// (21, 30, 'sp4_v_b_42')
// (21, 31, 'sp4_v_b_31')
// (21, 32, 'sp4_v_b_18')
// (21, 33, 'span4_horz_l_13')
// (21, 33, 'span4_vert_7')

reg io_26_33_0 = 0;
// (17, 20, 'neigh_op_tnr_5')
// (17, 21, 'neigh_op_rgt_5')
// (17, 21, 'sp12_h_r_1')
// (17, 22, 'neigh_op_bnr_5')
// (18, 20, 'neigh_op_top_5')
// (18, 21, 'lutff_5/out')
// (18, 21, 'sp12_h_r_2')
// (18, 22, 'neigh_op_bot_5')
// (19, 20, 'neigh_op_tnl_5')
// (19, 21, 'neigh_op_lft_5')
// (19, 21, 'sp12_h_r_5')
// (19, 22, 'neigh_op_bnl_5')
// (20, 21, 'sp12_h_r_6')
// (21, 21, 'sp12_h_r_9')
// (22, 21, 'sp12_h_r_10')
// (23, 21, 'sp12_h_r_13')
// (24, 21, 'sp12_h_r_14')
// (25, 21, 'sp12_h_r_17')
// (25, 33, 'span4_horz_r_3')
// (26, 21, 'sp12_h_r_18')
// (26, 33, 'io_0/D_OUT_0')
// (26, 33, 'io_0/PAD')
// (26, 33, 'local_g1_7')
// (26, 33, 'span4_horz_r_7')
// (27, 21, 'sp12_h_r_21')
// (27, 33, 'span4_horz_r_11')
// (28, 21, 'sp12_h_r_22')
// (28, 29, 'sp4_r_v_b_38')
// (28, 30, 'sp4_r_v_b_27')
// (28, 31, 'sp4_r_v_b_14')
// (28, 32, 'sp4_r_v_b_3')
// (28, 33, 'span4_horz_r_15')
// (29, 21, 'sp12_h_l_22')
// (29, 21, 'sp12_v_t_22')
// (29, 22, 'sp12_v_b_22')
// (29, 23, 'sp12_v_b_21')
// (29, 24, 'sp12_v_b_18')
// (29, 25, 'sp12_v_b_17')
// (29, 26, 'sp12_v_b_14')
// (29, 27, 'sp12_v_b_13')
// (29, 28, 'sp12_v_b_10')
// (29, 28, 'sp4_v_t_38')
// (29, 29, 'sp12_v_b_9')
// (29, 29, 'sp4_v_b_38')
// (29, 30, 'sp12_v_b_6')
// (29, 30, 'sp4_v_b_27')
// (29, 31, 'sp12_v_b_5')
// (29, 31, 'sp4_v_b_14')
// (29, 32, 'sp12_v_b_2')
// (29, 32, 'sp4_v_b_3')
// (29, 32, 'sp4_v_t_43')
// (29, 33, 'span12_vert_1')
// (29, 33, 'span4_horz_l_15')
// (29, 33, 'span4_vert_43')

reg io_20_33_0 = 0;
// (17, 20, 'neigh_op_tnr_7')
// (17, 21, 'neigh_op_rgt_7')
// (17, 22, 'neigh_op_bnr_7')
// (17, 26, 'sp4_r_v_b_36')
// (17, 27, 'sp4_r_v_b_25')
// (17, 28, 'sp4_r_v_b_12')
// (17, 29, 'sp4_r_v_b_1')
// (17, 30, 'sp4_r_v_b_36')
// (17, 31, 'sp4_r_v_b_25')
// (17, 32, 'sp4_r_v_b_12')
// (18, 16, 'sp12_v_t_22')
// (18, 17, 'sp12_v_b_22')
// (18, 18, 'sp12_v_b_21')
// (18, 19, 'sp12_v_b_18')
// (18, 20, 'neigh_op_top_7')
// (18, 20, 'sp12_v_b_17')
// (18, 21, 'lutff_7/out')
// (18, 21, 'sp12_v_b_14')
// (18, 22, 'neigh_op_bot_7')
// (18, 22, 'sp12_v_b_13')
// (18, 23, 'sp12_v_b_10')
// (18, 24, 'sp12_v_b_9')
// (18, 25, 'sp12_v_b_6')
// (18, 25, 'sp4_v_t_36')
// (18, 26, 'sp12_v_b_5')
// (18, 26, 'sp4_v_b_36')
// (18, 27, 'sp12_v_b_2')
// (18, 27, 'sp4_v_b_25')
// (18, 28, 'sp12_v_b_1')
// (18, 28, 'sp4_v_b_12')
// (18, 29, 'sp4_v_b_1')
// (18, 29, 'sp4_v_t_36')
// (18, 30, 'sp4_v_b_36')
// (18, 31, 'sp4_v_b_25')
// (18, 32, 'sp4_v_b_12')
// (18, 33, 'span4_horz_r_0')
// (18, 33, 'span4_vert_1')
// (19, 20, 'neigh_op_tnl_7')
// (19, 21, 'neigh_op_lft_7')
// (19, 22, 'neigh_op_bnl_7')
// (19, 33, 'span4_horz_r_4')
// (20, 33, 'io_0/D_OUT_0')
// (20, 33, 'io_0/PAD')
// (20, 33, 'local_g0_0')
// (20, 33, 'span4_horz_r_8')
// (21, 33, 'span4_horz_r_12')
// (22, 33, 'span4_horz_l_12')

reg n1256 = 0;
// (17, 20, 'sp4_r_v_b_43')
// (17, 21, 'sp4_r_v_b_30')
// (17, 22, 'sp4_r_v_b_19')
// (17, 23, 'sp4_r_v_b_6')
// (18, 19, 'sp4_h_r_0')
// (18, 19, 'sp4_v_t_43')
// (18, 20, 'local_g3_3')
// (18, 20, 'lutff_5/in_3')
// (18, 20, 'sp4_v_b_43')
// (18, 21, 'sp4_v_b_30')
// (18, 22, 'sp4_v_b_19')
// (18, 23, 'sp4_v_b_6')
// (19, 18, 'neigh_op_tnr_4')
// (19, 19, 'neigh_op_rgt_4')
// (19, 19, 'sp4_h_r_13')
// (19, 20, 'neigh_op_bnr_4')
// (20, 18, 'neigh_op_top_4')
// (20, 19, 'lutff_4/out')
// (20, 19, 'sp4_h_r_24')
// (20, 20, 'neigh_op_bot_4')
// (21, 18, 'neigh_op_tnl_4')
// (21, 19, 'neigh_op_lft_4')
// (21, 19, 'sp4_h_r_37')
// (21, 20, 'neigh_op_bnl_4')
// (22, 19, 'sp4_h_l_37')

reg n1257 = 0;
// (17, 21, 'local_g3_5')
// (17, 21, 'lutff_5/in_1')
// (17, 21, 'sp4_r_v_b_45')
// (17, 22, 'sp4_r_v_b_32')
// (17, 23, 'sp4_r_v_b_21')
// (17, 24, 'sp4_r_v_b_8')
// (18, 20, 'sp4_h_r_2')
// (18, 20, 'sp4_v_t_45')
// (18, 21, 'sp4_v_b_45')
// (18, 22, 'sp4_v_b_32')
// (18, 23, 'sp4_v_b_21')
// (18, 24, 'sp4_v_b_8')
// (19, 19, 'neigh_op_tnr_5')
// (19, 20, 'neigh_op_rgt_5')
// (19, 20, 'sp4_h_r_15')
// (19, 21, 'neigh_op_bnr_5')
// (20, 19, 'neigh_op_top_5')
// (20, 20, 'lutff_5/out')
// (20, 20, 'sp4_h_r_26')
// (20, 21, 'neigh_op_bot_5')
// (21, 19, 'neigh_op_tnl_5')
// (21, 20, 'neigh_op_lft_5')
// (21, 20, 'sp4_h_r_39')
// (21, 21, 'neigh_op_bnl_5')
// (22, 20, 'sp4_h_l_39')

wire n1258;
// (17, 21, 'neigh_op_tnr_3')
// (17, 22, 'neigh_op_rgt_3')
// (17, 23, 'neigh_op_bnr_3')
// (18, 21, 'neigh_op_top_3')
// (18, 22, 'lutff_3/out')
// (18, 23, 'neigh_op_bot_3')
// (19, 21, 'neigh_op_tnl_3')
// (19, 22, 'local_g0_3')
// (19, 22, 'local_g1_3')
// (19, 22, 'lutff_0/in_0')
// (19, 22, 'lutff_1/in_0')
// (19, 22, 'lutff_2/in_0')
// (19, 22, 'lutff_3/in_0')
// (19, 22, 'lutff_4/in_0')
// (19, 22, 'lutff_5/in_0')
// (19, 22, 'lutff_6/in_0')
// (19, 22, 'lutff_7/in_0')
// (19, 22, 'neigh_op_lft_3')
// (19, 23, 'neigh_op_bnl_3')

reg n1259 = 0;
// (17, 21, 'neigh_op_tnr_5')
// (17, 22, 'neigh_op_rgt_5')
// (17, 23, 'neigh_op_bnr_5')
// (18, 15, 'sp12_v_t_22')
// (18, 16, 'sp12_v_b_22')
// (18, 17, 'sp12_v_b_21')
// (18, 18, 'sp12_v_b_18')
// (18, 19, 'sp12_v_b_17')
// (18, 20, 'sp12_v_b_14')
// (18, 21, 'neigh_op_top_5')
// (18, 21, 'sp12_v_b_13')
// (18, 22, 'local_g3_5')
// (18, 22, 'lutff_5/in_1')
// (18, 22, 'lutff_5/out')
// (18, 22, 'sp12_v_b_10')
// (18, 23, 'neigh_op_bot_5')
// (18, 23, 'sp12_v_b_9')
// (18, 24, 'sp12_v_b_6')
// (18, 25, 'sp12_v_b_5')
// (18, 26, 'sp12_v_b_2')
// (18, 27, 'sp12_h_r_1')
// (18, 27, 'sp12_v_b_1')
// (19, 21, 'neigh_op_tnl_5')
// (19, 22, 'neigh_op_lft_5')
// (19, 23, 'neigh_op_bnl_5')
// (19, 27, 'sp12_h_r_2')
// (20, 27, 'sp12_h_r_5')
// (21, 27, 'sp12_h_r_6')
// (22, 27, 'sp12_h_r_9')
// (23, 27, 'sp12_h_r_10')
// (24, 27, 'sp12_h_r_13')
// (25, 27, 'sp12_h_r_14')
// (26, 27, 'sp12_h_r_17')
// (27, 27, 'sp12_h_r_18')
// (28, 27, 'sp12_h_r_21')
// (29, 27, 'sp12_h_r_22')
// (30, 15, 'sp12_h_r_1')
// (30, 15, 'sp12_v_t_22')
// (30, 16, 'sp12_v_b_22')
// (30, 17, 'sp12_v_b_21')
// (30, 18, 'sp12_v_b_18')
// (30, 19, 'sp12_v_b_17')
// (30, 20, 'sp12_v_b_14')
// (30, 21, 'sp12_v_b_13')
// (30, 22, 'sp12_v_b_10')
// (30, 23, 'sp12_v_b_9')
// (30, 24, 'sp12_v_b_6')
// (30, 25, 'sp12_v_b_5')
// (30, 26, 'sp12_v_b_2')
// (30, 27, 'sp12_h_l_22')
// (30, 27, 'sp12_v_b_1')
// (31, 15, 'sp12_h_r_2')
// (32, 15, 'sp12_h_r_5')
// (33, 15, 'io_0/OUT_ENB')
// (33, 15, 'local_g0_5')
// (33, 15, 'span12_horz_5')

reg n1260 = 0;
// (17, 21, 'neigh_op_tnr_6')
// (17, 22, 'neigh_op_rgt_6')
// (17, 23, 'neigh_op_bnr_6')
// (18, 16, 'sp12_h_r_0')
// (18, 16, 'sp12_v_t_23')
// (18, 17, 'sp12_v_b_23')
// (18, 18, 'sp12_v_b_20')
// (18, 19, 'sp12_v_b_19')
// (18, 20, 'sp12_v_b_16')
// (18, 21, 'neigh_op_top_6')
// (18, 21, 'sp12_v_b_15')
// (18, 22, 'local_g2_6')
// (18, 22, 'lutff_6/in_2')
// (18, 22, 'lutff_6/out')
// (18, 22, 'sp12_v_b_12')
// (18, 23, 'neigh_op_bot_6')
// (18, 23, 'sp12_v_b_11')
// (18, 24, 'sp12_v_b_8')
// (18, 25, 'sp12_v_b_7')
// (18, 26, 'sp12_v_b_4')
// (18, 27, 'sp12_v_b_3')
// (18, 28, 'sp12_v_b_0')
// (19, 16, 'sp12_h_r_3')
// (19, 21, 'neigh_op_tnl_6')
// (19, 22, 'neigh_op_lft_6')
// (19, 23, 'neigh_op_bnl_6')
// (20, 16, 'sp12_h_r_4')
// (21, 16, 'sp12_h_r_7')
// (22, 16, 'sp12_h_r_8')
// (23, 16, 'sp12_h_r_11')
// (24, 16, 'sp12_h_r_12')
// (25, 16, 'sp12_h_r_15')
// (26, 16, 'sp12_h_r_16')
// (27, 16, 'sp12_h_r_19')
// (28, 16, 'sp12_h_r_20')
// (29, 7, 'sp4_r_v_b_43')
// (29, 8, 'sp4_r_v_b_30')
// (29, 9, 'sp4_r_v_b_19')
// (29, 10, 'sp4_r_v_b_6')
// (29, 16, 'sp12_h_r_23')
// (30, 4, 'sp12_v_t_23')
// (30, 5, 'sp12_v_b_23')
// (30, 6, 'sp12_v_b_20')
// (30, 6, 'sp4_h_r_6')
// (30, 6, 'sp4_v_t_43')
// (30, 7, 'sp12_v_b_19')
// (30, 7, 'sp4_v_b_43')
// (30, 8, 'sp12_v_b_16')
// (30, 8, 'sp4_v_b_30')
// (30, 9, 'sp12_v_b_15')
// (30, 9, 'sp4_v_b_19')
// (30, 10, 'sp12_v_b_12')
// (30, 10, 'sp4_v_b_6')
// (30, 11, 'sp12_v_b_11')
// (30, 12, 'sp12_v_b_8')
// (30, 13, 'sp12_v_b_7')
// (30, 14, 'sp12_v_b_4')
// (30, 15, 'sp12_v_b_3')
// (30, 16, 'sp12_h_l_23')
// (30, 16, 'sp12_v_b_0')
// (31, 6, 'sp4_h_r_19')
// (32, 6, 'sp4_h_r_30')
// (33, 6, 'io_1/OUT_ENB')
// (33, 6, 'local_g0_6')
// (33, 6, 'span4_horz_30')

wire n1261;
// (17, 21, 'sp12_h_r_0')
// (18, 21, 'sp12_h_r_3')
// (19, 21, 'local_g0_4')
// (19, 21, 'lutff_2/in_2')
// (19, 21, 'sp12_h_r_4')
// (20, 21, 'sp12_h_r_7')
// (21, 21, 'sp12_h_r_8')
// (22, 21, 'sp12_h_r_11')
// (23, 21, 'sp12_h_r_12')
// (24, 21, 'sp12_h_r_15')
// (25, 21, 'sp12_h_r_16')
// (26, 21, 'sp12_h_r_19')
// (27, 21, 'sp12_h_r_20')
// (28, 21, 'sp12_h_r_23')
// (28, 32, 'neigh_op_tnr_0')
// (28, 32, 'neigh_op_tnr_4')
// (29, 21, 'sp12_h_l_23')
// (29, 21, 'sp12_v_t_23')
// (29, 22, 'sp12_v_b_23')
// (29, 23, 'sp12_v_b_20')
// (29, 24, 'sp12_v_b_19')
// (29, 25, 'sp12_v_b_16')
// (29, 26, 'sp12_v_b_15')
// (29, 27, 'sp12_v_b_12')
// (29, 28, 'sp12_v_b_11')
// (29, 29, 'sp12_v_b_8')
// (29, 30, 'sp12_v_b_7')
// (29, 31, 'sp12_v_b_4')
// (29, 32, 'neigh_op_top_0')
// (29, 32, 'neigh_op_top_4')
// (29, 32, 'sp12_v_b_3')
// (29, 33, 'io_0/D_IN_0')
// (29, 33, 'span12_vert_0')
// (30, 32, 'neigh_op_tnl_0')
// (30, 32, 'neigh_op_tnl_4')

reg n1262 = 0;
// (17, 21, 'sp4_r_v_b_44')
// (17, 22, 'sp4_r_v_b_33')
// (17, 23, 'sp4_r_v_b_20')
// (17, 24, 'sp4_r_v_b_9')
// (18, 20, 'sp4_h_r_3')
// (18, 20, 'sp4_v_t_44')
// (18, 21, 'sp4_v_b_44')
// (18, 22, 'sp4_v_b_33')
// (18, 23, 'sp4_v_b_20')
// (18, 24, 'local_g1_1')
// (18, 24, 'lutff_3/in_1')
// (18, 24, 'sp4_v_b_9')
// (19, 20, 'sp4_h_r_14')
// (20, 20, 'sp4_h_r_27')
// (21, 20, 'sp4_h_r_38')
// (22, 19, 'neigh_op_tnr_7')
// (22, 20, 'neigh_op_rgt_7')
// (22, 20, 'sp4_h_l_38')
// (22, 20, 'sp4_h_r_3')
// (22, 21, 'neigh_op_bnr_7')
// (23, 19, 'neigh_op_top_7')
// (23, 20, 'lutff_7/out')
// (23, 20, 'sp4_h_r_14')
// (23, 21, 'neigh_op_bot_7')
// (24, 19, 'neigh_op_tnl_7')
// (24, 20, 'neigh_op_lft_7')
// (24, 20, 'sp4_h_r_27')
// (24, 21, 'neigh_op_bnl_7')
// (25, 20, 'sp4_h_r_38')
// (26, 20, 'sp4_h_l_38')

wire n1263;
// (17, 22, 'lutff_7/cout')
// (17, 23, 'carry_in')
// (17, 23, 'carry_in_mux')

reg io_19_33_1 = 0;
// (17, 22, 'neigh_op_tnr_0')
// (17, 23, 'neigh_op_rgt_0')
// (17, 24, 'neigh_op_bnr_0')
// (18, 22, 'neigh_op_top_0')
// (18, 22, 'sp4_r_v_b_44')
// (18, 23, 'lutff_0/out')
// (18, 23, 'sp4_r_v_b_33')
// (18, 24, 'neigh_op_bot_0')
// (18, 24, 'sp4_r_v_b_20')
// (18, 25, 'sp4_r_v_b_9')
// (18, 26, 'sp4_r_v_b_44')
// (18, 27, 'sp4_r_v_b_33')
// (18, 28, 'sp4_r_v_b_20')
// (18, 29, 'sp4_r_v_b_9')
// (18, 30, 'sp4_r_v_b_44')
// (18, 31, 'sp4_r_v_b_33')
// (18, 32, 'sp4_r_v_b_20')
// (19, 21, 'sp4_v_t_44')
// (19, 22, 'neigh_op_tnl_0')
// (19, 22, 'sp4_v_b_44')
// (19, 23, 'neigh_op_lft_0')
// (19, 23, 'sp4_v_b_33')
// (19, 24, 'neigh_op_bnl_0')
// (19, 24, 'sp4_v_b_20')
// (19, 25, 'sp4_v_b_9')
// (19, 25, 'sp4_v_t_44')
// (19, 26, 'sp4_v_b_44')
// (19, 27, 'sp4_v_b_33')
// (19, 28, 'sp4_v_b_20')
// (19, 29, 'sp4_v_b_9')
// (19, 29, 'sp4_v_t_44')
// (19, 30, 'sp4_v_b_44')
// (19, 31, 'sp4_v_b_33')
// (19, 32, 'sp4_v_b_20')
// (19, 33, 'io_1/D_OUT_0')
// (19, 33, 'io_1/PAD')
// (19, 33, 'local_g0_1')
// (19, 33, 'span4_vert_9')

reg io_33_5_1 = 0;
// (17, 22, 'neigh_op_tnr_3')
// (17, 23, 'neigh_op_rgt_3')
// (17, 24, 'neigh_op_bnr_3')
// (18, 14, 'sp12_h_r_1')
// (18, 14, 'sp12_v_t_22')
// (18, 15, 'sp12_v_b_22')
// (18, 16, 'sp12_v_b_21')
// (18, 17, 'sp12_v_b_18')
// (18, 18, 'sp12_v_b_17')
// (18, 19, 'sp12_v_b_14')
// (18, 20, 'sp12_v_b_13')
// (18, 21, 'sp12_v_b_10')
// (18, 22, 'neigh_op_top_3')
// (18, 22, 'sp12_v_b_9')
// (18, 23, 'lutff_3/out')
// (18, 23, 'sp12_v_b_6')
// (18, 24, 'neigh_op_bot_3')
// (18, 24, 'sp12_v_b_5')
// (18, 25, 'sp12_v_b_2')
// (18, 26, 'sp12_v_b_1')
// (19, 14, 'sp12_h_r_2')
// (19, 22, 'neigh_op_tnl_3')
// (19, 23, 'neigh_op_lft_3')
// (19, 24, 'neigh_op_bnl_3')
// (20, 14, 'sp12_h_r_5')
// (21, 14, 'sp12_h_r_6')
// (22, 14, 'sp12_h_r_9')
// (23, 14, 'sp12_h_r_10')
// (24, 14, 'sp12_h_r_13')
// (25, 14, 'sp12_h_r_14')
// (26, 14, 'sp12_h_r_17')
// (27, 14, 'sp12_h_r_18')
// (28, 14, 'sp12_h_r_21')
// (29, 6, 'sp4_r_v_b_42')
// (29, 7, 'sp4_r_v_b_31')
// (29, 8, 'sp4_r_v_b_18')
// (29, 9, 'sp4_r_v_b_7')
// (29, 14, 'sp12_h_r_22')
// (30, 2, 'sp12_v_t_22')
// (30, 3, 'sp12_v_b_22')
// (30, 4, 'sp12_v_b_21')
// (30, 5, 'sp12_v_b_18')
// (30, 5, 'sp4_h_r_0')
// (30, 5, 'sp4_v_t_42')
// (30, 6, 'sp12_v_b_17')
// (30, 6, 'sp4_v_b_42')
// (30, 7, 'sp12_v_b_14')
// (30, 7, 'sp4_v_b_31')
// (30, 8, 'sp12_v_b_13')
// (30, 8, 'sp4_v_b_18')
// (30, 9, 'sp12_v_b_10')
// (30, 9, 'sp4_v_b_7')
// (30, 10, 'sp12_v_b_9')
// (30, 11, 'sp12_v_b_6')
// (30, 12, 'sp12_v_b_5')
// (30, 13, 'sp12_v_b_2')
// (30, 14, 'sp12_h_l_22')
// (30, 14, 'sp12_v_b_1')
// (31, 5, 'sp4_h_r_13')
// (32, 5, 'sp4_h_r_24')
// (33, 5, 'io_1/D_OUT_0')
// (33, 5, 'io_1/PAD')
// (33, 5, 'local_g1_0')
// (33, 5, 'span4_horz_24')

reg io_33_28_0 = 0;
// (17, 22, 'neigh_op_tnr_4')
// (17, 23, 'neigh_op_rgt_4')
// (17, 24, 'neigh_op_bnr_4')
// (18, 22, 'neigh_op_top_4')
// (18, 23, 'lutff_4/out')
// (18, 23, 'sp12_h_r_0')
// (18, 24, 'neigh_op_bot_4')
// (19, 22, 'neigh_op_tnl_4')
// (19, 23, 'neigh_op_lft_4')
// (19, 23, 'sp12_h_r_3')
// (19, 24, 'neigh_op_bnl_4')
// (20, 23, 'sp12_h_r_4')
// (21, 23, 'sp12_h_r_7')
// (22, 23, 'sp12_h_r_8')
// (23, 23, 'sp12_h_r_11')
// (24, 23, 'sp12_h_r_12')
// (25, 23, 'sp12_h_r_15')
// (25, 23, 'sp4_h_r_9')
// (26, 23, 'sp12_h_r_16')
// (26, 23, 'sp4_h_r_20')
// (27, 23, 'sp12_h_r_19')
// (27, 23, 'sp4_h_r_33')
// (28, 23, 'sp12_h_r_20')
// (28, 23, 'sp4_h_r_44')
// (29, 23, 'sp12_h_r_23')
// (29, 23, 'sp4_h_l_44')
// (29, 23, 'sp4_h_r_0')
// (30, 23, 'sp12_h_l_23')
// (30, 23, 'sp4_h_r_13')
// (31, 23, 'sp4_h_r_24')
// (32, 23, 'sp4_h_r_37')
// (33, 23, 'span4_horz_37')
// (33, 23, 'span4_vert_t_14')
// (33, 24, 'span4_vert_b_14')
// (33, 25, 'span4_vert_b_10')
// (33, 26, 'span4_vert_b_6')
// (33, 27, 'span4_vert_b_2')
// (33, 27, 'span4_vert_t_14')
// (33, 28, 'io_0/D_OUT_0')
// (33, 28, 'io_0/PAD')
// (33, 28, 'local_g0_6')
// (33, 28, 'span4_vert_b_14')
// (33, 29, 'span4_vert_b_10')
// (33, 30, 'span4_vert_b_6')
// (33, 31, 'span4_vert_b_2')

reg io_25_33_0 = 0;
// (17, 22, 'neigh_op_tnr_5')
// (17, 23, 'neigh_op_rgt_5')
// (17, 23, 'sp4_r_v_b_42')
// (17, 24, 'neigh_op_bnr_5')
// (17, 24, 'sp4_r_v_b_31')
// (17, 25, 'sp4_r_v_b_18')
// (17, 26, 'sp4_r_v_b_7')
// (17, 27, 'sp4_r_v_b_42')
// (17, 28, 'sp4_r_v_b_31')
// (17, 29, 'sp4_r_v_b_18')
// (17, 30, 'sp4_r_v_b_7')
// (18, 22, 'neigh_op_top_5')
// (18, 22, 'sp4_v_t_42')
// (18, 23, 'lutff_5/out')
// (18, 23, 'sp4_v_b_42')
// (18, 24, 'neigh_op_bot_5')
// (18, 24, 'sp4_v_b_31')
// (18, 25, 'sp4_v_b_18')
// (18, 26, 'sp4_v_b_7')
// (18, 26, 'sp4_v_t_42')
// (18, 27, 'sp4_v_b_42')
// (18, 28, 'sp4_v_b_31')
// (18, 29, 'sp4_v_b_18')
// (18, 30, 'sp4_h_r_7')
// (18, 30, 'sp4_v_b_7')
// (19, 22, 'neigh_op_tnl_5')
// (19, 23, 'neigh_op_lft_5')
// (19, 24, 'neigh_op_bnl_5')
// (19, 30, 'sp4_h_r_18')
// (20, 30, 'sp4_h_r_31')
// (21, 30, 'sp4_h_r_42')
// (21, 31, 'sp4_r_v_b_37')
// (21, 32, 'sp4_r_v_b_24')
// (22, 30, 'sp4_h_l_42')
// (22, 30, 'sp4_v_t_37')
// (22, 31, 'sp4_v_b_37')
// (22, 32, 'sp4_v_b_24')
// (22, 33, 'span4_horz_r_2')
// (22, 33, 'span4_vert_13')
// (23, 33, 'span4_horz_r_6')
// (24, 33, 'span4_horz_r_10')
// (25, 33, 'io_0/D_OUT_0')
// (25, 33, 'io_0/PAD')
// (25, 33, 'local_g0_6')
// (25, 33, 'span4_horz_r_14')
// (26, 33, 'span4_horz_l_14')

reg io_33_21_0 = 0;
// (17, 22, 'neigh_op_tnr_7')
// (17, 23, 'neigh_op_rgt_7')
// (17, 23, 'sp4_h_r_3')
// (17, 24, 'neigh_op_bnr_7')
// (18, 22, 'neigh_op_top_7')
// (18, 23, 'lutff_7/out')
// (18, 23, 'sp4_h_r_14')
// (18, 24, 'neigh_op_bot_7')
// (19, 22, 'neigh_op_tnl_7')
// (19, 23, 'neigh_op_lft_7')
// (19, 23, 'sp4_h_r_27')
// (19, 24, 'neigh_op_bnl_7')
// (20, 23, 'sp4_h_r_38')
// (21, 23, 'sp4_h_l_38')
// (21, 23, 'sp4_h_r_3')
// (22, 23, 'sp4_h_r_14')
// (23, 23, 'sp4_h_r_27')
// (24, 23, 'sp4_h_r_38')
// (25, 23, 'sp4_h_l_38')
// (25, 23, 'sp4_h_r_6')
// (26, 23, 'sp4_h_r_19')
// (27, 23, 'sp4_h_r_30')
// (28, 23, 'sp4_h_r_43')
// (29, 23, 'sp4_h_l_43')
// (29, 23, 'sp4_h_r_6')
// (30, 23, 'sp4_h_r_19')
// (31, 23, 'sp4_h_r_30')
// (32, 23, 'sp4_h_r_43')
// (33, 19, 'span4_vert_t_15')
// (33, 20, 'span4_vert_b_15')
// (33, 21, 'io_0/D_OUT_0')
// (33, 21, 'io_0/PAD')
// (33, 21, 'local_g1_3')
// (33, 21, 'span4_vert_b_11')
// (33, 22, 'span4_vert_b_7')
// (33, 23, 'span4_horz_43')
// (33, 23, 'span4_vert_b_3')

wire n1269;
// (17, 23, 'lutff_7/cout')
// (17, 24, 'carry_in')
// (17, 24, 'carry_in_mux')

wire n1270;
// (17, 23, 'neigh_op_tnr_1')
// (17, 24, 'neigh_op_rgt_1')
// (17, 25, 'neigh_op_bnr_1')
// (18, 23, 'neigh_op_top_1')
// (18, 24, 'local_g2_1')
// (18, 24, 'lutff_1/out')
// (18, 24, 'lutff_4/in_3')
// (18, 25, 'neigh_op_bot_1')
// (19, 23, 'neigh_op_tnl_1')
// (19, 24, 'neigh_op_lft_1')
// (19, 25, 'neigh_op_bnl_1')

wire n1271;
// (17, 23, 'neigh_op_tnr_2')
// (17, 24, 'neigh_op_rgt_2')
// (17, 25, 'neigh_op_bnr_2')
// (18, 23, 'neigh_op_top_2')
// (18, 24, 'local_g2_2')
// (18, 24, 'lutff_2/out')
// (18, 24, 'lutff_5/in_3')
// (18, 25, 'neigh_op_bot_2')
// (19, 23, 'neigh_op_tnl_2')
// (19, 24, 'neigh_op_lft_2')
// (19, 25, 'neigh_op_bnl_2')

reg n1272 = 0;
// (17, 23, 'neigh_op_tnr_6')
// (17, 24, 'neigh_op_rgt_6')
// (17, 25, 'neigh_op_bnr_6')
// (18, 23, 'neigh_op_top_6')
// (18, 24, 'local_g0_6')
// (18, 24, 'lutff_3/in_3')
// (18, 24, 'lutff_6/out')
// (18, 25, 'neigh_op_bot_6')
// (19, 23, 'neigh_op_tnl_6')
// (19, 24, 'neigh_op_lft_6')
// (19, 25, 'neigh_op_bnl_6')

reg n1273 = 0;
// (17, 23, 'sp4_r_v_b_39')
// (17, 24, 'sp4_r_v_b_26')
// (17, 25, 'sp4_r_v_b_15')
// (17, 26, 'sp4_r_v_b_2')
// (18, 22, 'local_g0_2')
// (18, 22, 'local_g1_2')
// (18, 22, 'lutff_3/in_0')
// (18, 22, 'lutff_4/in_2')
// (18, 22, 'sp4_h_r_2')
// (18, 22, 'sp4_v_t_39')
// (18, 23, 'sp4_v_b_39')
// (18, 24, 'sp4_v_b_26')
// (18, 25, 'sp4_v_b_15')
// (18, 26, 'local_g0_2')
// (18, 26, 'lutff_0/in_2')
// (18, 26, 'sp4_v_b_2')
// (19, 21, 'neigh_op_tnr_5')
// (19, 22, 'neigh_op_rgt_5')
// (19, 22, 'sp4_h_r_15')
// (19, 23, 'neigh_op_bnr_5')
// (20, 21, 'neigh_op_top_5')
// (20, 22, 'local_g2_5')
// (20, 22, 'lutff_1/in_0')
// (20, 22, 'lutff_5/in_2')
// (20, 22, 'lutff_5/out')
// (20, 22, 'sp4_h_r_26')
// (20, 23, 'neigh_op_bot_5')
// (21, 21, 'neigh_op_tnl_5')
// (21, 22, 'neigh_op_lft_5')
// (21, 22, 'sp4_h_r_39')
// (21, 23, 'neigh_op_bnl_5')
// (22, 22, 'sp4_h_l_39')

wire n1274;
// (17, 24, 'lutff_7/cout')
// (17, 25, 'carry_in')
// (17, 25, 'carry_in_mux')
// (17, 25, 'lutff_0/in_3')

wire n1275;
// (17, 24, 'neigh_op_tnr_2')
// (17, 25, 'neigh_op_rgt_2')
// (17, 26, 'neigh_op_bnr_2')
// (18, 15, 'sp12_v_t_23')
// (18, 16, 'sp12_v_b_23')
// (18, 17, 'sp12_v_b_20')
// (18, 18, 'sp12_v_b_19')
// (18, 19, 'sp12_v_b_16')
// (18, 20, 'local_g3_7')
// (18, 20, 'lutff_7/in_1')
// (18, 20, 'sp12_v_b_15')
// (18, 21, 'sp12_v_b_12')
// (18, 22, 'sp12_v_b_11')
// (18, 23, 'sp12_v_b_8')
// (18, 24, 'neigh_op_top_2')
// (18, 24, 'sp12_v_b_7')
// (18, 25, 'lutff_2/out')
// (18, 25, 'sp12_v_b_4')
// (18, 26, 'neigh_op_bot_2')
// (18, 26, 'sp12_v_b_3')
// (18, 27, 'sp12_v_b_0')
// (19, 24, 'neigh_op_tnl_2')
// (19, 25, 'neigh_op_lft_2')
// (19, 26, 'neigh_op_bnl_2')

wire n1276;
// (17, 24, 'neigh_op_tnr_3')
// (17, 25, 'neigh_op_rgt_3')
// (17, 26, 'neigh_op_bnr_3')
// (18, 24, 'local_g1_3')
// (18, 24, 'lutff_7/in_1')
// (18, 24, 'neigh_op_top_3')
// (18, 25, 'lutff_3/out')
// (18, 26, 'neigh_op_bot_3')
// (19, 24, 'neigh_op_tnl_3')
// (19, 25, 'neigh_op_lft_3')
// (19, 26, 'neigh_op_bnl_3')

wire n1277;
// (17, 24, 'neigh_op_tnr_4')
// (17, 25, 'neigh_op_rgt_4')
// (17, 26, 'neigh_op_bnr_4')
// (18, 24, 'local_g0_4')
// (18, 24, 'lutff_5/in_1')
// (18, 24, 'neigh_op_top_4')
// (18, 25, 'lutff_4/out')
// (18, 26, 'neigh_op_bot_4')
// (19, 24, 'neigh_op_tnl_4')
// (19, 25, 'neigh_op_lft_4')
// (19, 26, 'neigh_op_bnl_4')

wire n1278;
// (17, 24, 'neigh_op_tnr_5')
// (17, 25, 'neigh_op_rgt_5')
// (17, 26, 'neigh_op_bnr_5')
// (18, 24, 'local_g1_5')
// (18, 24, 'lutff_7/in_3')
// (18, 24, 'neigh_op_top_5')
// (18, 25, 'lutff_5/out')
// (18, 26, 'neigh_op_bot_5')
// (19, 24, 'neigh_op_tnl_5')
// (19, 25, 'neigh_op_lft_5')
// (19, 26, 'neigh_op_bnl_5')

wire n1279;
// (17, 24, 'neigh_op_tnr_6')
// (17, 25, 'neigh_op_rgt_6')
// (17, 25, 'sp4_r_v_b_44')
// (17, 26, 'neigh_op_bnr_6')
// (17, 26, 'sp4_r_v_b_33')
// (17, 27, 'sp4_r_v_b_20')
// (17, 28, 'sp4_r_v_b_9')
// (18, 24, 'neigh_op_top_6')
// (18, 24, 'sp4_h_r_9')
// (18, 24, 'sp4_v_t_44')
// (18, 25, 'lutff_6/out')
// (18, 25, 'sp4_v_b_44')
// (18, 26, 'neigh_op_bot_6')
// (18, 26, 'sp4_v_b_33')
// (18, 27, 'sp4_v_b_20')
// (18, 28, 'sp4_v_b_9')
// (19, 24, 'neigh_op_tnl_6')
// (19, 24, 'sp4_h_r_20')
// (19, 25, 'neigh_op_lft_6')
// (19, 26, 'neigh_op_bnl_6')
// (20, 24, 'sp4_h_r_33')
// (21, 21, 'local_g2_6')
// (21, 21, 'lutff_1/in_3')
// (21, 21, 'sp4_r_v_b_38')
// (21, 22, 'sp4_r_v_b_27')
// (21, 23, 'sp4_r_v_b_14')
// (21, 24, 'sp4_h_r_44')
// (21, 24, 'sp4_r_v_b_3')
// (22, 20, 'sp4_v_t_38')
// (22, 21, 'sp4_v_b_38')
// (22, 22, 'sp4_v_b_27')
// (22, 23, 'sp4_v_b_14')
// (22, 24, 'sp4_h_l_44')
// (22, 24, 'sp4_v_b_3')

wire n1280;
// (17, 25, 'neigh_op_tnr_5')
// (17, 26, 'neigh_op_rgt_5')
// (17, 27, 'neigh_op_bnr_5')
// (18, 19, 'sp12_v_t_22')
// (18, 20, 'local_g2_6')
// (18, 20, 'lutff_1/in_3')
// (18, 20, 'sp12_v_b_22')
// (18, 21, 'sp12_v_b_21')
// (18, 22, 'sp12_v_b_18')
// (18, 23, 'sp12_v_b_17')
// (18, 24, 'sp12_v_b_14')
// (18, 25, 'neigh_op_top_5')
// (18, 25, 'sp12_v_b_13')
// (18, 26, 'lutff_5/out')
// (18, 26, 'sp12_v_b_10')
// (18, 27, 'neigh_op_bot_5')
// (18, 27, 'sp12_v_b_9')
// (18, 28, 'sp12_v_b_6')
// (18, 29, 'sp12_v_b_5')
// (18, 30, 'sp12_v_b_2')
// (18, 31, 'sp12_v_b_1')
// (19, 25, 'neigh_op_tnl_5')
// (19, 26, 'neigh_op_lft_5')
// (19, 27, 'neigh_op_bnl_5')

reg n1281 = 0;
// (17, 25, 'sp4_h_r_3')
// (18, 25, 'local_g0_6')
// (18, 25, 'lutff_5/in_1')
// (18, 25, 'sp4_h_r_14')
// (19, 19, 'neigh_op_tnr_7')
// (19, 20, 'neigh_op_rgt_7')
// (19, 21, 'neigh_op_bnr_7')
// (19, 25, 'sp4_h_r_27')
// (20, 18, 'sp4_r_v_b_39')
// (20, 19, 'neigh_op_top_7')
// (20, 19, 'sp4_r_v_b_26')
// (20, 20, 'lutff_7/out')
// (20, 20, 'sp4_r_v_b_15')
// (20, 21, 'neigh_op_bot_7')
// (20, 21, 'sp4_r_v_b_2')
// (20, 22, 'sp4_r_v_b_47')
// (20, 23, 'sp4_r_v_b_34')
// (20, 24, 'sp4_r_v_b_23')
// (20, 25, 'sp4_h_r_38')
// (20, 25, 'sp4_r_v_b_10')
// (21, 17, 'sp4_v_t_39')
// (21, 18, 'sp4_v_b_39')
// (21, 19, 'neigh_op_tnl_7')
// (21, 19, 'sp4_v_b_26')
// (21, 20, 'neigh_op_lft_7')
// (21, 20, 'sp4_v_b_15')
// (21, 21, 'neigh_op_bnl_7')
// (21, 21, 'sp4_v_b_2')
// (21, 21, 'sp4_v_t_47')
// (21, 22, 'sp4_v_b_47')
// (21, 23, 'sp4_v_b_34')
// (21, 24, 'sp4_v_b_23')
// (21, 25, 'sp4_h_l_38')
// (21, 25, 'sp4_v_b_10')

reg n1282 = 0;
// (17, 26, 'sp4_h_r_6')
// (18, 26, 'local_g1_3')
// (18, 26, 'lutff_5/in_1')
// (18, 26, 'sp4_h_r_19')
// (19, 26, 'sp4_h_r_30')
// (20, 22, 'neigh_op_tnr_2')
// (20, 23, 'neigh_op_rgt_2')
// (20, 23, 'sp4_r_v_b_36')
// (20, 24, 'neigh_op_bnr_2')
// (20, 24, 'sp4_r_v_b_25')
// (20, 25, 'sp4_r_v_b_12')
// (20, 26, 'sp4_h_r_43')
// (20, 26, 'sp4_r_v_b_1')
// (21, 22, 'neigh_op_top_2')
// (21, 22, 'sp4_v_t_36')
// (21, 23, 'lutff_2/out')
// (21, 23, 'sp4_v_b_36')
// (21, 24, 'neigh_op_bot_2')
// (21, 24, 'sp4_v_b_25')
// (21, 25, 'sp4_v_b_12')
// (21, 26, 'sp4_h_l_43')
// (21, 26, 'sp4_v_b_1')
// (22, 22, 'neigh_op_tnl_2')
// (22, 23, 'neigh_op_lft_2')
// (22, 24, 'neigh_op_bnl_2')

reg n1283 = 0;
// (18, 0, 'span12_vert_17')
// (18, 1, 'sp12_v_b_17')
// (18, 2, 'sp12_v_b_14')
// (18, 3, 'sp12_v_b_13')
// (18, 4, 'sp12_v_b_10')
// (18, 5, 'sp12_v_b_9')
// (18, 6, 'sp12_v_b_6')
// (18, 7, 'sp12_v_b_5')
// (18, 8, 'sp12_v_b_2')
// (18, 9, 'local_g3_1')
// (18, 9, 'lutff_5/in_3')
// (18, 9, 'sp12_v_b_1')
// (18, 9, 'sp12_v_t_22')
// (18, 10, 'sp12_v_b_22')
// (18, 11, 'sp12_v_b_21')
// (18, 12, 'sp12_v_b_18')
// (18, 13, 'sp12_v_b_17')
// (18, 14, 'sp12_v_b_14')
// (18, 15, 'sp12_v_b_13')
// (18, 16, 'sp12_v_b_10')
// (18, 17, 'sp12_v_b_9')
// (18, 18, 'sp12_v_b_6')
// (18, 19, 'sp12_v_b_5')
// (18, 20, 'neigh_op_tnr_5')
// (18, 20, 'sp12_v_b_2')
// (18, 21, 'neigh_op_rgt_5')
// (18, 21, 'sp12_h_r_1')
// (18, 21, 'sp12_v_b_1')
// (18, 22, 'neigh_op_bnr_5')
// (19, 20, 'neigh_op_top_5')
// (19, 21, 'lutff_5/out')
// (19, 21, 'sp12_h_r_2')
// (19, 22, 'neigh_op_bot_5')
// (20, 20, 'neigh_op_tnl_5')
// (20, 21, 'neigh_op_lft_5')
// (20, 21, 'sp12_h_r_5')
// (20, 22, 'neigh_op_bnl_5')
// (21, 21, 'sp12_h_r_6')
// (22, 21, 'sp12_h_r_9')
// (23, 21, 'sp12_h_r_10')
// (24, 21, 'sp12_h_r_13')
// (25, 21, 'sp12_h_r_14')
// (26, 21, 'sp12_h_r_17')
// (27, 21, 'sp12_h_r_18')
// (28, 21, 'sp12_h_r_21')
// (29, 21, 'sp12_h_r_22')
// (30, 21, 'sp12_h_l_22')

reg n1284 = 0;
// (18, 8, 'sp4_r_v_b_39')
// (18, 9, 'local_g0_2')
// (18, 9, 'lutff_3/in_3')
// (18, 9, 'sp4_r_v_b_26')
// (18, 10, 'sp4_r_v_b_15')
// (18, 11, 'sp4_r_v_b_2')
// (18, 12, 'sp4_r_v_b_46')
// (18, 13, 'sp4_r_v_b_35')
// (18, 14, 'sp4_r_v_b_22')
// (18, 15, 'sp4_r_v_b_11')
// (18, 20, 'neigh_op_tnr_3')
// (18, 21, 'neigh_op_rgt_3')
// (18, 22, 'neigh_op_bnr_3')
// (19, 7, 'sp4_v_t_39')
// (19, 8, 'sp4_v_b_39')
// (19, 9, 'sp4_v_b_26')
// (19, 10, 'sp4_v_b_15')
// (19, 11, 'sp4_v_b_2')
// (19, 11, 'sp4_v_t_46')
// (19, 12, 'sp12_v_t_22')
// (19, 12, 'sp4_v_b_46')
// (19, 13, 'sp12_v_b_22')
// (19, 13, 'sp4_v_b_35')
// (19, 14, 'sp12_v_b_21')
// (19, 14, 'sp4_v_b_22')
// (19, 15, 'sp12_v_b_18')
// (19, 15, 'sp4_v_b_11')
// (19, 16, 'sp12_v_b_17')
// (19, 17, 'sp12_v_b_14')
// (19, 18, 'sp12_v_b_13')
// (19, 19, 'sp12_v_b_10')
// (19, 20, 'neigh_op_top_3')
// (19, 20, 'sp12_v_b_9')
// (19, 21, 'lutff_3/out')
// (19, 21, 'sp12_v_b_6')
// (19, 22, 'neigh_op_bot_3')
// (19, 22, 'sp12_v_b_5')
// (19, 23, 'sp12_v_b_2')
// (19, 24, 'sp12_v_b_1')
// (20, 20, 'neigh_op_tnl_3')
// (20, 21, 'neigh_op_lft_3')
// (20, 22, 'neigh_op_bnl_3')

reg n1285 = 0;
// (18, 8, 'sp4_r_v_b_41')
// (18, 9, 'local_g1_4')
// (18, 9, 'lutff_6/in_3')
// (18, 9, 'sp4_r_v_b_28')
// (18, 10, 'sp4_r_v_b_17')
// (18, 11, 'sp4_r_v_b_4')
// (18, 20, 'neigh_op_tnr_6')
// (18, 21, 'neigh_op_rgt_6')
// (18, 22, 'neigh_op_bnr_6')
// (19, 3, 'sp12_v_t_23')
// (19, 4, 'sp12_v_b_23')
// (19, 5, 'sp12_v_b_20')
// (19, 6, 'sp12_v_b_19')
// (19, 7, 'sp12_v_b_16')
// (19, 7, 'sp4_v_t_41')
// (19, 8, 'sp12_v_b_15')
// (19, 8, 'sp4_v_b_41')
// (19, 9, 'sp12_v_b_12')
// (19, 9, 'sp4_v_b_28')
// (19, 10, 'sp12_v_b_11')
// (19, 10, 'sp4_v_b_17')
// (19, 11, 'sp12_v_b_8')
// (19, 11, 'sp4_v_b_4')
// (19, 12, 'sp12_v_b_7')
// (19, 13, 'sp12_v_b_4')
// (19, 14, 'sp12_v_b_3')
// (19, 15, 'sp12_v_b_0')
// (19, 15, 'sp12_v_t_23')
// (19, 16, 'sp12_v_b_23')
// (19, 17, 'sp12_v_b_20')
// (19, 18, 'sp12_v_b_19')
// (19, 19, 'sp12_v_b_16')
// (19, 20, 'neigh_op_top_6')
// (19, 20, 'sp12_v_b_15')
// (19, 21, 'lutff_6/out')
// (19, 21, 'sp12_v_b_12')
// (19, 22, 'neigh_op_bot_6')
// (19, 22, 'sp12_v_b_11')
// (19, 23, 'sp12_v_b_8')
// (19, 24, 'sp12_v_b_7')
// (19, 25, 'sp12_v_b_4')
// (19, 26, 'sp12_v_b_3')
// (19, 27, 'sp12_v_b_0')
// (20, 20, 'neigh_op_tnl_6')
// (20, 21, 'neigh_op_lft_6')
// (20, 22, 'neigh_op_bnl_6')

reg n1286 = 0;
// (18, 8, 'sp4_r_v_b_42')
// (18, 9, 'local_g1_7')
// (18, 9, 'lutff_7/in_3')
// (18, 9, 'sp4_r_v_b_31')
// (18, 10, 'sp4_r_v_b_18')
// (18, 11, 'sp4_r_v_b_7')
// (18, 20, 'neigh_op_tnr_7')
// (18, 21, 'neigh_op_rgt_7')
// (18, 22, 'neigh_op_bnr_7')
// (19, 4, 'sp12_v_t_22')
// (19, 5, 'sp12_v_b_22')
// (19, 6, 'sp12_v_b_21')
// (19, 7, 'sp12_v_b_18')
// (19, 7, 'sp4_v_t_42')
// (19, 8, 'sp12_v_b_17')
// (19, 8, 'sp4_v_b_42')
// (19, 9, 'sp12_v_b_14')
// (19, 9, 'sp4_v_b_31')
// (19, 10, 'sp12_v_b_13')
// (19, 10, 'sp4_v_b_18')
// (19, 11, 'sp12_v_b_10')
// (19, 11, 'sp4_v_b_7')
// (19, 12, 'sp12_v_b_9')
// (19, 13, 'sp12_v_b_6')
// (19, 14, 'sp12_v_b_5')
// (19, 15, 'sp12_v_b_2')
// (19, 16, 'sp12_v_b_1')
// (19, 16, 'sp12_v_t_22')
// (19, 17, 'sp12_v_b_22')
// (19, 18, 'sp12_v_b_21')
// (19, 19, 'sp12_v_b_18')
// (19, 20, 'neigh_op_top_7')
// (19, 20, 'sp12_v_b_17')
// (19, 21, 'lutff_7/out')
// (19, 21, 'sp12_v_b_14')
// (19, 22, 'neigh_op_bot_7')
// (19, 22, 'sp12_v_b_13')
// (19, 23, 'sp12_v_b_10')
// (19, 24, 'sp12_v_b_9')
// (19, 25, 'sp12_v_b_6')
// (19, 26, 'sp12_v_b_5')
// (19, 27, 'sp12_v_b_2')
// (19, 28, 'sp12_v_b_1')
// (20, 20, 'neigh_op_tnl_7')
// (20, 21, 'neigh_op_lft_7')
// (20, 22, 'neigh_op_bnl_7')

reg n1287 = 0;
// (18, 8, 'sp4_r_v_b_43')
// (18, 9, 'local_g1_6')
// (18, 9, 'lutff_4/in_3')
// (18, 9, 'sp4_r_v_b_30')
// (18, 10, 'sp4_r_v_b_19')
// (18, 11, 'sp4_r_v_b_6')
// (18, 12, 'sp4_r_v_b_47')
// (18, 13, 'sp4_r_v_b_34')
// (18, 14, 'sp4_r_v_b_23')
// (18, 15, 'sp4_r_v_b_10')
// (18, 20, 'neigh_op_tnr_4')
// (18, 21, 'neigh_op_rgt_4')
// (18, 22, 'neigh_op_bnr_4')
// (19, 7, 'sp4_v_t_43')
// (19, 8, 'sp4_v_b_43')
// (19, 9, 'sp4_v_b_30')
// (19, 10, 'sp4_v_b_19')
// (19, 11, 'sp4_v_b_6')
// (19, 11, 'sp4_v_t_47')
// (19, 12, 'sp4_v_b_47')
// (19, 13, 'sp12_v_t_23')
// (19, 13, 'sp4_v_b_34')
// (19, 14, 'sp12_v_b_23')
// (19, 14, 'sp4_v_b_23')
// (19, 15, 'sp12_v_b_20')
// (19, 15, 'sp4_v_b_10')
// (19, 16, 'sp12_v_b_19')
// (19, 17, 'sp12_v_b_16')
// (19, 18, 'sp12_v_b_15')
// (19, 19, 'sp12_v_b_12')
// (19, 20, 'neigh_op_top_4')
// (19, 20, 'sp12_v_b_11')
// (19, 21, 'lutff_4/out')
// (19, 21, 'sp12_v_b_8')
// (19, 22, 'neigh_op_bot_4')
// (19, 22, 'sp12_v_b_7')
// (19, 23, 'sp12_v_b_4')
// (19, 24, 'sp12_v_b_3')
// (19, 25, 'sp12_v_b_0')
// (20, 20, 'neigh_op_tnl_4')
// (20, 21, 'neigh_op_lft_4')
// (20, 22, 'neigh_op_bnl_4')

reg n1288 = 0;
// (18, 8, 'sp4_r_v_b_45')
// (18, 9, 'local_g0_3')
// (18, 9, 'lutff_2/in_3')
// (18, 9, 'sp4_r_v_b_32')
// (18, 10, 'sp4_r_v_b_21')
// (18, 11, 'sp4_r_v_b_8')
// (18, 20, 'neigh_op_tnr_2')
// (18, 21, 'neigh_op_rgt_2')
// (18, 22, 'neigh_op_bnr_2')
// (19, 7, 'sp12_v_t_23')
// (19, 7, 'sp4_v_t_45')
// (19, 8, 'sp12_v_b_23')
// (19, 8, 'sp4_v_b_45')
// (19, 9, 'sp12_v_b_20')
// (19, 9, 'sp4_v_b_32')
// (19, 10, 'sp12_v_b_19')
// (19, 10, 'sp4_v_b_21')
// (19, 11, 'sp12_v_b_16')
// (19, 11, 'sp4_v_b_8')
// (19, 12, 'sp12_v_b_15')
// (19, 13, 'sp12_v_b_12')
// (19, 14, 'sp12_v_b_11')
// (19, 15, 'sp12_v_b_8')
// (19, 16, 'sp12_v_b_7')
// (19, 17, 'sp12_v_b_4')
// (19, 18, 'sp12_v_b_3')
// (19, 19, 'sp12_v_b_0')
// (19, 19, 'sp12_v_t_23')
// (19, 20, 'neigh_op_top_2')
// (19, 20, 'sp12_v_b_23')
// (19, 21, 'lutff_2/out')
// (19, 21, 'sp12_v_b_20')
// (19, 22, 'neigh_op_bot_2')
// (19, 22, 'sp12_v_b_19')
// (19, 23, 'sp12_v_b_16')
// (19, 24, 'sp12_v_b_15')
// (19, 25, 'sp12_v_b_12')
// (19, 26, 'sp12_v_b_11')
// (19, 27, 'sp12_v_b_8')
// (19, 28, 'sp12_v_b_7')
// (19, 29, 'sp12_v_b_4')
// (19, 30, 'sp12_v_b_3')
// (19, 31, 'sp12_v_b_0')
// (20, 20, 'neigh_op_tnl_2')
// (20, 21, 'neigh_op_lft_2')
// (20, 22, 'neigh_op_bnl_2')

reg n1289 = 0;
// (18, 9, 'neigh_op_tnr_0')
// (18, 10, 'neigh_op_rgt_0')
// (18, 11, 'neigh_op_bnr_0')
// (19, 6, 'sp12_v_t_23')
// (19, 7, 'sp12_v_b_23')
// (19, 8, 'sp12_v_b_20')
// (19, 9, 'neigh_op_top_0')
// (19, 9, 'sp12_v_b_19')
// (19, 10, 'lutff_0/out')
// (19, 10, 'sp12_v_b_16')
// (19, 11, 'neigh_op_bot_0')
// (19, 11, 'sp12_v_b_15')
// (19, 12, 'sp12_v_b_12')
// (19, 13, 'local_g3_3')
// (19, 13, 'lutff_5/in_1')
// (19, 13, 'sp12_v_b_11')
// (19, 14, 'sp12_v_b_8')
// (19, 15, 'sp12_v_b_7')
// (19, 16, 'sp12_v_b_4')
// (19, 17, 'sp12_v_b_3')
// (19, 18, 'sp12_v_b_0')
// (20, 9, 'neigh_op_tnl_0')
// (20, 10, 'neigh_op_lft_0')
// (20, 11, 'neigh_op_bnl_0')

reg n1290 = 0;
// (18, 9, 'neigh_op_tnr_2')
// (18, 10, 'neigh_op_rgt_2')
// (18, 10, 'sp4_h_r_9')
// (18, 11, 'neigh_op_bnr_2')
// (19, 9, 'neigh_op_top_2')
// (19, 10, 'lutff_2/out')
// (19, 10, 'sp4_h_r_20')
// (19, 11, 'neigh_op_bot_2')
// (20, 9, 'neigh_op_tnl_2')
// (20, 10, 'neigh_op_lft_2')
// (20, 10, 'sp4_h_r_33')
// (20, 11, 'neigh_op_bnl_2')
// (21, 10, 'sp4_h_r_44')
// (21, 11, 'sp4_r_v_b_39')
// (21, 12, 'sp4_r_v_b_26')
// (21, 13, 'sp4_r_v_b_15')
// (21, 14, 'sp4_r_v_b_2')
// (21, 15, 'sp4_r_v_b_39')
// (21, 16, 'local_g0_2')
// (21, 16, 'lutff_1/in_1')
// (21, 16, 'sp4_r_v_b_26')
// (21, 17, 'sp4_r_v_b_15')
// (21, 18, 'sp4_r_v_b_2')
// (22, 10, 'sp4_h_l_44')
// (22, 10, 'sp4_v_t_39')
// (22, 11, 'sp4_v_b_39')
// (22, 12, 'sp4_v_b_26')
// (22, 13, 'sp4_v_b_15')
// (22, 14, 'sp4_v_b_2')
// (22, 14, 'sp4_v_t_39')
// (22, 15, 'sp4_v_b_39')
// (22, 16, 'sp4_v_b_26')
// (22, 17, 'sp4_v_b_15')
// (22, 18, 'sp4_v_b_2')

reg n1291 = 0;
// (18, 9, 'neigh_op_tnr_4')
// (18, 10, 'neigh_op_rgt_4')
// (18, 11, 'neigh_op_bnr_4')
// (19, 9, 'neigh_op_top_4')
// (19, 10, 'lutff_4/out')
// (19, 10, 'sp12_h_r_0')
// (19, 10, 'sp12_v_t_23')
// (19, 11, 'neigh_op_bot_4')
// (19, 11, 'sp12_v_b_23')
// (19, 12, 'sp12_v_b_20')
// (19, 13, 'sp12_v_b_19')
// (19, 14, 'sp12_v_b_16')
// (19, 15, 'sp12_v_b_15')
// (19, 16, 'sp12_v_b_12')
// (19, 17, 'sp12_v_b_11')
// (19, 18, 'local_g2_0')
// (19, 18, 'lutff_1/in_1')
// (19, 18, 'sp12_v_b_8')
// (19, 19, 'sp12_v_b_7')
// (19, 20, 'sp12_v_b_4')
// (19, 21, 'sp12_v_b_3')
// (19, 22, 'sp12_v_b_0')
// (20, 9, 'neigh_op_tnl_4')
// (20, 10, 'neigh_op_lft_4')
// (20, 10, 'sp12_h_r_3')
// (20, 11, 'neigh_op_bnl_4')
// (21, 10, 'sp12_h_r_4')
// (22, 10, 'sp12_h_r_7')
// (23, 10, 'sp12_h_r_8')
// (24, 10, 'sp12_h_r_11')
// (25, 10, 'sp12_h_r_12')
// (26, 10, 'sp12_h_r_15')
// (27, 10, 'sp12_h_r_16')
// (28, 10, 'sp12_h_r_19')
// (29, 10, 'sp12_h_r_20')
// (30, 10, 'sp12_h_r_23')
// (31, 10, 'sp12_h_l_23')

reg n1292 = 0;
// (18, 9, 'neigh_op_tnr_5')
// (18, 10, 'neigh_op_rgt_5')
// (18, 11, 'neigh_op_bnr_5')
// (19, 3, 'sp12_v_t_22')
// (19, 4, 'sp12_v_b_22')
// (19, 5, 'sp12_v_b_21')
// (19, 6, 'sp12_v_b_18')
// (19, 7, 'sp12_v_b_17')
// (19, 8, 'sp12_v_b_14')
// (19, 9, 'neigh_op_top_5')
// (19, 9, 'sp12_v_b_13')
// (19, 10, 'lutff_5/out')
// (19, 10, 'sp12_v_b_10')
// (19, 11, 'neigh_op_bot_5')
// (19, 11, 'sp12_v_b_9')
// (19, 12, 'sp12_v_b_6')
// (19, 13, 'sp12_v_b_5')
// (19, 14, 'local_g2_2')
// (19, 14, 'lutff_1/in_1')
// (19, 14, 'sp12_v_b_2')
// (19, 15, 'sp12_v_b_1')
// (20, 9, 'neigh_op_tnl_5')
// (20, 10, 'neigh_op_lft_5')
// (20, 11, 'neigh_op_bnl_5')

wire n1293;
// (18, 9, 'sp12_v_t_23')
// (18, 10, 'sp12_v_b_23')
// (18, 11, 'sp12_v_b_20')
// (18, 12, 'sp12_v_b_19')
// (18, 13, 'local_g3_0')
// (18, 13, 'lutff_2/in_3')
// (18, 13, 'sp12_v_b_16')
// (18, 14, 'sp12_v_b_15')
// (18, 15, 'sp12_v_b_12')
// (18, 16, 'sp12_v_b_11')
// (18, 17, 'sp12_v_b_8')
// (18, 18, 'sp12_v_b_7')
// (18, 19, 'sp12_v_b_4')
// (18, 20, 'sp12_v_b_3')
// (18, 21, 'sp12_h_r_0')
// (18, 21, 'sp12_v_b_0')
// (19, 20, 'neigh_op_tnr_6')
// (19, 21, 'neigh_op_rgt_6')
// (19, 21, 'sp12_h_r_3')
// (19, 22, 'neigh_op_bnr_6')
// (20, 20, 'neigh_op_top_6')
// (20, 21, 'lutff_6/out')
// (20, 21, 'sp12_h_r_4')
// (20, 22, 'neigh_op_bot_6')
// (21, 20, 'neigh_op_tnl_6')
// (21, 21, 'neigh_op_lft_6')
// (21, 21, 'sp12_h_r_7')
// (21, 22, 'neigh_op_bnl_6')
// (22, 21, 'sp12_h_r_8')
// (23, 21, 'sp12_h_r_11')
// (24, 21, 'sp12_h_r_12')
// (25, 21, 'sp12_h_r_15')
// (26, 21, 'sp12_h_r_16')
// (27, 21, 'sp12_h_r_19')
// (28, 21, 'sp12_h_r_20')
// (29, 21, 'sp12_h_r_23')
// (30, 21, 'sp12_h_l_23')

reg n1294 = 0;
// (18, 9, 'sp4_h_r_11')
// (19, 9, 'sp4_h_r_22')
// (20, 9, 'local_g3_3')
// (20, 9, 'lutff_7/in_1')
// (20, 9, 'sp4_h_r_35')
// (21, 9, 'neigh_op_tnr_4')
// (21, 9, 'sp4_h_r_46')
// (21, 10, 'local_g3_4')
// (21, 10, 'lutff_4/in_1')
// (21, 10, 'lutff_7/in_0')
// (21, 10, 'neigh_op_rgt_4')
// (21, 10, 'sp4_r_v_b_40')
// (21, 11, 'neigh_op_bnr_4')
// (21, 11, 'sp4_r_v_b_29')
// (21, 12, 'sp4_r_v_b_16')
// (21, 13, 'sp4_r_v_b_5')
// (22, 9, 'neigh_op_top_4')
// (22, 9, 'sp4_h_l_46')
// (22, 9, 'sp4_v_t_40')
// (22, 10, 'local_g3_4')
// (22, 10, 'lutff_4/in_1')
// (22, 10, 'lutff_4/out')
// (22, 10, 'sp4_v_b_40')
// (22, 11, 'neigh_op_bot_4')
// (22, 11, 'sp4_v_b_29')
// (22, 12, 'sp4_v_b_16')
// (22, 13, 'sp4_v_b_5')
// (23, 9, 'neigh_op_tnl_4')
// (23, 10, 'neigh_op_lft_4')
// (23, 11, 'neigh_op_bnl_4')

reg n1295 = 0;
// (18, 10, 'neigh_op_tnr_1')
// (18, 11, 'neigh_op_rgt_1')
// (18, 12, 'neigh_op_bnr_1')
// (19, 10, 'neigh_op_top_1')
// (19, 10, 'sp4_r_v_b_46')
// (19, 11, 'lutff_1/out')
// (19, 11, 'sp4_r_v_b_35')
// (19, 12, 'neigh_op_bot_1')
// (19, 12, 'sp4_r_v_b_22')
// (19, 13, 'sp4_r_v_b_11')
// (20, 9, 'sp4_v_t_46')
// (20, 10, 'neigh_op_tnl_1')
// (20, 10, 'sp4_v_b_46')
// (20, 11, 'neigh_op_lft_1')
// (20, 11, 'sp4_v_b_35')
// (20, 12, 'neigh_op_bnl_1')
// (20, 12, 'sp4_v_b_22')
// (20, 13, 'local_g0_3')
// (20, 13, 'lutff_0/in_3')
// (20, 13, 'sp4_v_b_11')

reg n1296 = 0;
// (18, 10, 'neigh_op_tnr_2')
// (18, 11, 'neigh_op_rgt_2')
// (18, 12, 'neigh_op_bnr_2')
// (19, 10, 'neigh_op_top_2')
// (19, 11, 'lutff_2/out')
// (19, 11, 'sp4_r_v_b_37')
// (19, 12, 'neigh_op_bot_2')
// (19, 12, 'sp4_r_v_b_24')
// (19, 13, 'sp4_r_v_b_13')
// (19, 14, 'sp4_r_v_b_0')
// (20, 10, 'neigh_op_tnl_2')
// (20, 10, 'sp4_v_t_37')
// (20, 11, 'neigh_op_lft_2')
// (20, 11, 'sp4_v_b_37')
// (20, 12, 'neigh_op_bnl_2')
// (20, 12, 'sp4_v_b_24')
// (20, 13, 'local_g0_5')
// (20, 13, 'lutff_6/in_3')
// (20, 13, 'sp4_v_b_13')
// (20, 14, 'sp4_v_b_0')

reg n1297 = 0;
// (18, 10, 'neigh_op_tnr_3')
// (18, 11, 'neigh_op_rgt_3')
// (18, 11, 'sp4_h_r_11')
// (18, 12, 'neigh_op_bnr_3')
// (19, 10, 'neigh_op_top_3')
// (19, 11, 'lutff_3/out')
// (19, 11, 'sp4_h_r_22')
// (19, 12, 'neigh_op_bot_3')
// (20, 10, 'neigh_op_tnl_3')
// (20, 11, 'neigh_op_lft_3')
// (20, 11, 'sp4_h_r_35')
// (20, 12, 'neigh_op_bnl_3')
// (21, 11, 'sp4_h_r_46')
// (21, 12, 'sp4_r_v_b_41')
// (21, 13, 'sp4_r_v_b_28')
// (21, 14, 'sp4_r_v_b_17')
// (21, 15, 'local_g1_4')
// (21, 15, 'lutff_0/in_3')
// (21, 15, 'sp4_r_v_b_4')
// (22, 11, 'sp4_h_l_46')
// (22, 11, 'sp4_v_t_41')
// (22, 12, 'sp4_v_b_41')
// (22, 13, 'sp4_v_b_28')
// (22, 14, 'sp4_v_b_17')
// (22, 15, 'sp4_v_b_4')

wire n1298;
// (18, 11, 'neigh_op_tnr_1')
// (18, 11, 'sp4_r_v_b_47')
// (18, 12, 'local_g2_2')
// (18, 12, 'lutff_global/cen')
// (18, 12, 'neigh_op_rgt_1')
// (18, 12, 'sp4_r_v_b_34')
// (18, 13, 'neigh_op_bnr_1')
// (18, 13, 'sp4_r_v_b_23')
// (18, 14, 'sp4_r_v_b_10')
// (19, 10, 'sp4_v_t_47')
// (19, 11, 'neigh_op_top_1')
// (19, 11, 'sp4_v_b_47')
// (19, 12, 'lutff_1/out')
// (19, 12, 'sp4_v_b_34')
// (19, 13, 'neigh_op_bot_1')
// (19, 13, 'sp4_v_b_23')
// (19, 14, 'sp4_v_b_10')
// (20, 11, 'neigh_op_tnl_1')
// (20, 12, 'neigh_op_lft_1')
// (20, 13, 'neigh_op_bnl_1')

wire n1299;
// (18, 11, 'neigh_op_tnr_2')
// (18, 12, 'neigh_op_rgt_2')
// (18, 13, 'neigh_op_bnr_2')
// (19, 11, 'neigh_op_top_2')
// (19, 12, 'lutff_2/out')
// (19, 13, 'neigh_op_bot_2')
// (20, 11, 'neigh_op_tnl_2')
// (20, 12, 'local_g0_2')
// (20, 12, 'lutff_global/cen')
// (20, 12, 'neigh_op_lft_2')
// (20, 13, 'neigh_op_bnl_2')

wire n1300;
// (18, 11, 'neigh_op_tnr_3')
// (18, 12, 'neigh_op_rgt_3')
// (18, 13, 'neigh_op_bnr_3')
// (19, 11, 'local_g1_3')
// (19, 11, 'lutff_global/cen')
// (19, 11, 'neigh_op_top_3')
// (19, 12, 'lutff_3/out')
// (19, 13, 'neigh_op_bot_3')
// (20, 11, 'neigh_op_tnl_3')
// (20, 12, 'neigh_op_lft_3')
// (20, 13, 'neigh_op_bnl_3')

wire n1301;
// (18, 11, 'neigh_op_tnr_4')
// (18, 12, 'neigh_op_rgt_4')
// (18, 13, 'neigh_op_bnr_4')
// (19, 11, 'neigh_op_top_4')
// (19, 12, 'lutff_4/out')
// (19, 12, 'sp4_h_r_8')
// (19, 13, 'neigh_op_bot_4')
// (20, 11, 'neigh_op_tnl_4')
// (20, 12, 'neigh_op_lft_4')
// (20, 12, 'sp4_h_r_21')
// (20, 13, 'neigh_op_bnl_4')
// (21, 12, 'sp4_h_r_32')
// (22, 12, 'sp4_h_r_45')
// (23, 12, 'local_g1_3')
// (23, 12, 'lutff_global/cen')
// (23, 12, 'sp4_h_l_45')
// (23, 12, 'sp4_h_r_11')
// (24, 12, 'sp4_h_r_22')
// (25, 12, 'sp4_h_r_35')
// (26, 12, 'sp4_h_r_46')
// (27, 12, 'sp4_h_l_46')

wire n1302;
// (18, 11, 'neigh_op_tnr_6')
// (18, 12, 'neigh_op_rgt_6')
// (18, 13, 'neigh_op_bnr_6')
// (19, 11, 'neigh_op_top_6')
// (19, 12, 'local_g2_6')
// (19, 12, 'lutff_5/in_3')
// (19, 12, 'lutff_6/out')
// (19, 12, 'sp4_r_v_b_45')
// (19, 13, 'neigh_op_bot_6')
// (19, 13, 'sp4_r_v_b_32')
// (19, 14, 'sp4_r_v_b_21')
// (19, 15, 'sp4_r_v_b_8')
// (20, 11, 'neigh_op_tnl_6')
// (20, 11, 'sp4_v_t_45')
// (20, 12, 'neigh_op_lft_6')
// (20, 12, 'sp4_v_b_45')
// (20, 13, 'neigh_op_bnl_6')
// (20, 13, 'sp4_v_b_32')
// (20, 14, 'sp4_v_b_21')
// (20, 15, 'local_g1_0')
// (20, 15, 'lutff_3/in_0')
// (20, 15, 'lutff_4/in_3')
// (20, 15, 'lutff_6/in_3')
// (20, 15, 'sp4_v_b_8')

reg n1303 = 0;
// (18, 12, 'neigh_op_tnr_0')
// (18, 13, 'neigh_op_rgt_0')
// (18, 14, 'neigh_op_bnr_0')
// (19, 12, 'neigh_op_top_0')
// (19, 13, 'local_g1_0')
// (19, 13, 'lutff_0/out')
// (19, 13, 'lutff_6/in_3')
// (19, 14, 'neigh_op_bot_0')
// (20, 12, 'neigh_op_tnl_0')
// (20, 13, 'neigh_op_lft_0')
// (20, 14, 'neigh_op_bnl_0')

wire n1304;
// (18, 12, 'neigh_op_tnr_3')
// (18, 13, 'neigh_op_rgt_3')
// (18, 14, 'neigh_op_bnr_3')
// (19, 12, 'neigh_op_top_3')
// (19, 13, 'lutff_3/out')
// (19, 14, 'neigh_op_bot_3')
// (20, 12, 'neigh_op_tnl_3')
// (20, 13, 'neigh_op_lft_3')
// (20, 14, 'local_g3_3')
// (20, 14, 'lutff_1/in_1')
// (20, 14, 'neigh_op_bnl_3')

wire n1305;
// (18, 12, 'neigh_op_tnr_4')
// (18, 13, 'neigh_op_rgt_4')
// (18, 14, 'neigh_op_bnr_4')
// (19, 12, 'neigh_op_top_4')
// (19, 13, 'local_g0_4')
// (19, 13, 'lutff_3/in_3')
// (19, 13, 'lutff_4/out')
// (19, 14, 'neigh_op_bot_4')
// (20, 12, 'neigh_op_tnl_4')
// (20, 13, 'neigh_op_lft_4')
// (20, 14, 'neigh_op_bnl_4')

wire n1306;
// (18, 12, 'neigh_op_tnr_6')
// (18, 13, 'neigh_op_rgt_6')
// (18, 14, 'local_g1_6')
// (18, 14, 'lutff_2/in_1')
// (18, 14, 'neigh_op_bnr_6')
// (19, 12, 'neigh_op_top_6')
// (19, 13, 'lutff_6/out')
// (19, 14, 'neigh_op_bot_6')
// (20, 12, 'neigh_op_tnl_6')
// (20, 13, 'neigh_op_lft_6')
// (20, 14, 'neigh_op_bnl_6')

wire n1307;
// (18, 12, 'neigh_op_tnr_7')
// (18, 13, 'neigh_op_rgt_7')
// (18, 14, 'neigh_op_bnr_7')
// (19, 12, 'neigh_op_top_7')
// (19, 13, 'local_g2_7')
// (19, 13, 'lutff_4/in_3')
// (19, 13, 'lutff_7/out')
// (19, 14, 'neigh_op_bot_7')
// (20, 12, 'neigh_op_tnl_7')
// (20, 13, 'neigh_op_lft_7')
// (20, 14, 'neigh_op_bnl_7')

reg n1308 = 0;
// (18, 12, 'sp4_h_r_0')
// (19, 11, 'neigh_op_tnr_4')
// (19, 12, 'neigh_op_rgt_4')
// (19, 12, 'sp4_h_r_13')
// (19, 13, 'neigh_op_bnr_4')
// (20, 11, 'neigh_op_top_4')
// (20, 12, 'lutff_4/out')
// (20, 12, 'sp4_h_r_24')
// (20, 13, 'neigh_op_bot_4')
// (21, 11, 'neigh_op_tnl_4')
// (21, 12, 'neigh_op_lft_4')
// (21, 12, 'sp4_h_r_37')
// (21, 13, 'neigh_op_bnl_4')
// (21, 13, 'sp4_r_v_b_37')
// (21, 14, 'sp4_r_v_b_24')
// (21, 15, 'sp4_r_v_b_13')
// (21, 16, 'sp4_r_v_b_0')
// (22, 12, 'sp4_h_l_37')
// (22, 12, 'sp4_v_t_37')
// (22, 13, 'local_g2_5')
// (22, 13, 'lutff_4/in_3')
// (22, 13, 'sp4_v_b_37')
// (22, 14, 'sp4_v_b_24')
// (22, 15, 'sp4_v_b_13')
// (22, 16, 'sp4_v_b_0')

reg n1309 = 0;
// (18, 12, 'sp4_h_r_2')
// (19, 11, 'neigh_op_tnr_5')
// (19, 12, 'neigh_op_rgt_5')
// (19, 12, 'sp4_h_r_15')
// (19, 13, 'neigh_op_bnr_5')
// (20, 11, 'neigh_op_top_5')
// (20, 12, 'lutff_5/out')
// (20, 12, 'sp4_h_r_26')
// (20, 13, 'neigh_op_bot_5')
// (21, 11, 'neigh_op_tnl_5')
// (21, 12, 'neigh_op_lft_5')
// (21, 12, 'sp4_h_r_39')
// (21, 13, 'neigh_op_bnl_5')
// (21, 13, 'sp4_r_v_b_39')
// (21, 14, 'sp4_r_v_b_26')
// (21, 15, 'sp4_r_v_b_15')
// (21, 16, 'sp4_r_v_b_2')
// (22, 12, 'sp4_h_l_39')
// (22, 12, 'sp4_v_t_39')
// (22, 13, 'local_g3_7')
// (22, 13, 'lutff_7/in_3')
// (22, 13, 'sp4_v_b_39')
// (22, 14, 'sp4_v_b_26')
// (22, 15, 'sp4_v_b_15')
// (22, 16, 'sp4_v_b_2')

wire n1310;
// (18, 13, 'local_g0_0')
// (18, 13, 'lutff_3/in_1')
// (18, 13, 'sp4_h_r_8')
// (19, 13, 'sp4_h_r_21')
// (20, 13, 'sp4_h_r_32')
// (21, 13, 'sp4_h_r_45')
// (21, 14, 'sp4_r_v_b_45')
// (21, 15, 'sp4_r_v_b_32')
// (21, 16, 'sp4_r_v_b_21')
// (21, 17, 'sp4_r_v_b_8')
// (21, 18, 'neigh_op_tnr_4')
// (21, 18, 'sp4_r_v_b_37')
// (21, 19, 'neigh_op_rgt_4')
// (21, 19, 'sp4_r_v_b_24')
// (21, 20, 'neigh_op_bnr_4')
// (21, 20, 'sp4_r_v_b_13')
// (21, 21, 'sp4_r_v_b_0')
// (22, 13, 'sp4_h_l_45')
// (22, 13, 'sp4_v_t_45')
// (22, 14, 'sp4_v_b_45')
// (22, 15, 'sp4_v_b_32')
// (22, 16, 'sp4_v_b_21')
// (22, 17, 'sp4_v_b_8')
// (22, 17, 'sp4_v_t_37')
// (22, 18, 'neigh_op_top_4')
// (22, 18, 'sp4_v_b_37')
// (22, 19, 'lutff_4/out')
// (22, 19, 'sp4_v_b_24')
// (22, 20, 'neigh_op_bot_4')
// (22, 20, 'sp4_v_b_13')
// (22, 21, 'sp4_v_b_0')
// (23, 18, 'neigh_op_tnl_4')
// (23, 19, 'neigh_op_lft_4')
// (23, 20, 'neigh_op_bnl_4')

wire n1311;
// (18, 13, 'local_g3_5')
// (18, 13, 'lutff_0/in_0')
// (18, 13, 'neigh_op_tnr_5')
// (18, 14, 'neigh_op_rgt_5')
// (18, 15, 'neigh_op_bnr_5')
// (19, 13, 'neigh_op_top_5')
// (19, 14, 'lutff_5/out')
// (19, 15, 'neigh_op_bot_5')
// (20, 13, 'neigh_op_tnl_5')
// (20, 14, 'neigh_op_lft_5')
// (20, 15, 'neigh_op_bnl_5')

wire n1312;
// (18, 13, 'lutff_0/lout')
// (18, 13, 'lutff_1/in_2')

wire n1313;
// (18, 13, 'lutff_2/lout')
// (18, 13, 'lutff_3/in_2')

wire n1314;
// (18, 13, 'lutff_3/lout')
// (18, 13, 'lutff_4/in_2')

wire n1315;
// (18, 13, 'lutff_6/lout')
// (18, 13, 'lutff_7/in_2')

reg n1316 = 0;
// (18, 13, 'neigh_op_tnr_0')
// (18, 14, 'neigh_op_rgt_0')
// (18, 15, 'neigh_op_bnr_0')
// (19, 13, 'neigh_op_top_0')
// (19, 14, 'local_g1_0')
// (19, 14, 'lutff_0/out')
// (19, 14, 'lutff_2/in_3')
// (19, 15, 'neigh_op_bot_0')
// (20, 13, 'neigh_op_tnl_0')
// (20, 14, 'neigh_op_lft_0')
// (20, 15, 'neigh_op_bnl_0')

wire n1317;
// (18, 13, 'neigh_op_tnr_2')
// (18, 14, 'neigh_op_rgt_2')
// (18, 14, 'sp4_r_v_b_36')
// (18, 15, 'neigh_op_bnr_2')
// (18, 15, 'sp4_r_v_b_25')
// (18, 16, 'sp4_r_v_b_12')
// (18, 17, 'sp4_r_v_b_1')
// (19, 13, 'neigh_op_top_2')
// (19, 13, 'sp4_v_t_36')
// (19, 14, 'lutff_2/out')
// (19, 14, 'sp4_v_b_36')
// (19, 15, 'neigh_op_bot_2')
// (19, 15, 'sp4_v_b_25')
// (19, 16, 'sp4_v_b_12')
// (19, 17, 'local_g1_1')
// (19, 17, 'lutff_3/in_1')
// (19, 17, 'sp4_v_b_1')
// (20, 13, 'neigh_op_tnl_2')
// (20, 14, 'neigh_op_lft_2')
// (20, 15, 'neigh_op_bnl_2')

wire n1318;
// (18, 13, 'neigh_op_tnr_6')
// (18, 14, 'neigh_op_rgt_6')
// (18, 15, 'neigh_op_bnr_6')
// (19, 13, 'neigh_op_top_6')
// (19, 14, 'local_g2_6')
// (19, 14, 'lutff_5/in_3')
// (19, 14, 'lutff_6/out')
// (19, 15, 'neigh_op_bot_6')
// (20, 13, 'neigh_op_tnl_6')
// (20, 14, 'neigh_op_lft_6')
// (20, 15, 'neigh_op_bnl_6')

wire n1319;
// (18, 13, 'neigh_op_tnr_7')
// (18, 14, 'neigh_op_rgt_7')
// (18, 15, 'neigh_op_bnr_7')
// (19, 13, 'neigh_op_top_7')
// (19, 14, 'local_g2_7')
// (19, 14, 'lutff_6/in_3')
// (19, 14, 'lutff_7/out')
// (19, 15, 'neigh_op_bot_7')
// (20, 13, 'neigh_op_tnl_7')
// (20, 14, 'neigh_op_lft_7')
// (20, 15, 'neigh_op_bnl_7')

reg n1320 = 0;
// (18, 13, 'sp12_v_t_23')
// (18, 14, 'sp12_v_b_23')
// (18, 15, 'sp12_v_b_20')
// (18, 16, 'sp12_v_b_19')
// (18, 17, 'sp12_v_b_16')
// (18, 18, 'local_g2_7')
// (18, 18, 'lutff_4/in_1')
// (18, 18, 'sp12_v_b_15')
// (18, 19, 'sp12_v_b_12')
// (18, 20, 'sp12_v_b_11')
// (18, 21, 'sp12_v_b_8')
// (18, 22, 'sp12_v_b_7')
// (18, 23, 'sp12_v_b_4')
// (18, 24, 'sp12_v_b_3')
// (18, 25, 'sp12_h_r_0')
// (18, 25, 'sp12_v_b_0')
// (19, 24, 'neigh_op_tnr_6')
// (19, 25, 'neigh_op_rgt_6')
// (19, 25, 'sp12_h_r_3')
// (19, 26, 'neigh_op_bnr_6')
// (20, 24, 'neigh_op_top_6')
// (20, 25, 'lutff_6/out')
// (20, 25, 'sp12_h_r_4')
// (20, 26, 'neigh_op_bot_6')
// (21, 24, 'neigh_op_tnl_6')
// (21, 25, 'neigh_op_lft_6')
// (21, 25, 'sp12_h_r_7')
// (21, 26, 'neigh_op_bnl_6')
// (22, 25, 'sp12_h_r_8')
// (23, 25, 'sp12_h_r_11')
// (24, 25, 'sp12_h_r_12')
// (25, 25, 'sp12_h_r_15')
// (26, 25, 'sp12_h_r_16')
// (27, 25, 'sp12_h_r_19')
// (28, 25, 'sp12_h_r_20')
// (29, 25, 'sp12_h_r_23')
// (30, 25, 'sp12_h_l_23')

reg n1321 = 0;
// (18, 13, 'sp4_r_v_b_39')
// (18, 14, 'sp4_r_v_b_26')
// (18, 15, 'neigh_op_tnr_1')
// (18, 15, 'sp4_r_v_b_15')
// (18, 16, 'neigh_op_rgt_1')
// (18, 16, 'sp4_r_v_b_2')
// (18, 17, 'neigh_op_bnr_1')
// (19, 12, 'sp4_v_t_39')
// (19, 13, 'local_g3_7')
// (19, 13, 'lutff_7/in_1')
// (19, 13, 'sp4_v_b_39')
// (19, 14, 'sp4_v_b_26')
// (19, 15, 'neigh_op_top_1')
// (19, 15, 'sp4_v_b_15')
// (19, 16, 'lutff_1/out')
// (19, 16, 'sp4_v_b_2')
// (19, 17, 'neigh_op_bot_1')
// (20, 15, 'neigh_op_tnl_1')
// (20, 16, 'neigh_op_lft_1')
// (20, 17, 'neigh_op_bnl_1')

reg n1322 = 0;
// (18, 13, 'sp4_r_v_b_43')
// (18, 14, 'sp4_r_v_b_30')
// (18, 15, 'sp4_r_v_b_19')
// (18, 16, 'sp4_r_v_b_6')
// (19, 12, 'sp4_v_t_43')
// (19, 13, 'sp4_v_b_43')
// (19, 14, 'sp4_v_b_30')
// (19, 15, 'local_g1_3')
// (19, 15, 'lutff_7/in_3')
// (19, 15, 'sp4_v_b_19')
// (19, 16, 'sp4_h_r_1')
// (19, 16, 'sp4_v_b_6')
// (20, 16, 'sp4_h_r_12')
// (21, 16, 'sp4_h_r_25')
// (22, 16, 'sp4_h_r_36')
// (23, 15, 'neigh_op_tnr_0')
// (23, 16, 'neigh_op_rgt_0')
// (23, 16, 'sp4_h_l_36')
// (23, 16, 'sp4_h_r_5')
// (23, 17, 'neigh_op_bnr_0')
// (24, 15, 'neigh_op_top_0')
// (24, 16, 'lutff_0/out')
// (24, 16, 'sp4_h_r_16')
// (24, 17, 'neigh_op_bot_0')
// (25, 15, 'neigh_op_tnl_0')
// (25, 16, 'neigh_op_lft_0')
// (25, 16, 'sp4_h_r_29')
// (25, 17, 'neigh_op_bnl_0')
// (26, 16, 'sp4_h_r_40')
// (27, 16, 'sp4_h_l_40')

wire n1323;
// (18, 14, 'local_g3_2')
// (18, 14, 'lutff_2/in_3')
// (18, 14, 'neigh_op_tnr_2')
// (18, 15, 'neigh_op_rgt_2')
// (18, 16, 'neigh_op_bnr_2')
// (19, 14, 'neigh_op_top_2')
// (19, 15, 'lutff_2/out')
// (19, 16, 'neigh_op_bot_2')
// (20, 14, 'neigh_op_tnl_2')
// (20, 15, 'neigh_op_lft_2')
// (20, 16, 'neigh_op_bnl_2')

wire n1324;
// (18, 14, 'lutff_0/lout')
// (18, 14, 'lutff_1/in_2')

wire n1325;
// (18, 14, 'lutff_2/lout')
// (18, 14, 'lutff_3/in_2')

wire n1326;
// (18, 14, 'lutff_4/lout')
// (18, 14, 'lutff_5/in_2')

reg n1327 = 0;
// (18, 14, 'neigh_op_tnr_0')
// (18, 15, 'neigh_op_rgt_0')
// (18, 16, 'neigh_op_bnr_0')
// (19, 14, 'neigh_op_top_0')
// (19, 15, 'local_g1_0')
// (19, 15, 'lutff_0/out')
// (19, 15, 'lutff_2/in_3')
// (19, 16, 'neigh_op_bot_0')
// (20, 14, 'neigh_op_tnl_0')
// (20, 15, 'neigh_op_lft_0')
// (20, 16, 'neigh_op_bnl_0')

wire n1328;
// (18, 14, 'neigh_op_tnr_4')
// (18, 15, 'neigh_op_rgt_4')
// (18, 16, 'neigh_op_bnr_4')
// (19, 14, 'neigh_op_top_4')
// (19, 15, 'lutff_4/out')
// (19, 16, 'neigh_op_bot_4')
// (20, 14, 'local_g3_4')
// (20, 14, 'lutff_6/in_1')
// (20, 14, 'neigh_op_tnl_4')
// (20, 15, 'neigh_op_lft_4')
// (20, 16, 'neigh_op_bnl_4')

reg n1329 = 0;
// (18, 14, 'neigh_op_tnr_5')
// (18, 15, 'neigh_op_rgt_5')
// (18, 16, 'neigh_op_bnr_5')
// (19, 14, 'neigh_op_top_5')
// (19, 15, 'local_g2_5')
// (19, 15, 'lutff_4/in_3')
// (19, 15, 'lutff_5/out')
// (19, 16, 'neigh_op_bot_5')
// (20, 14, 'neigh_op_tnl_5')
// (20, 15, 'neigh_op_lft_5')
// (20, 16, 'neigh_op_bnl_5')

wire n1330;
// (18, 14, 'neigh_op_tnr_7')
// (18, 15, 'neigh_op_rgt_7')
// (18, 15, 'sp4_h_r_3')
// (18, 16, 'neigh_op_bnr_7')
// (19, 14, 'neigh_op_top_7')
// (19, 15, 'lutff_7/out')
// (19, 15, 'sp4_h_r_14')
// (19, 16, 'neigh_op_bot_7')
// (20, 14, 'neigh_op_tnl_7')
// (20, 15, 'neigh_op_lft_7')
// (20, 15, 'sp4_h_r_27')
// (20, 16, 'neigh_op_bnl_7')
// (21, 15, 'sp4_h_r_38')
// (21, 16, 'sp4_r_v_b_38')
// (21, 17, 'sp4_r_v_b_27')
// (21, 18, 'sp4_r_v_b_14')
// (21, 19, 'local_g1_3')
// (21, 19, 'lutff_3/in_3')
// (21, 19, 'sp4_r_v_b_3')
// (22, 15, 'sp4_h_l_38')
// (22, 15, 'sp4_v_t_38')
// (22, 16, 'sp4_v_b_38')
// (22, 17, 'sp4_v_b_27')
// (22, 18, 'sp4_v_b_14')
// (22, 19, 'sp4_v_b_3')

reg n1331 = 0;
// (18, 14, 'sp4_r_v_b_44')
// (18, 15, 'neigh_op_tnr_2')
// (18, 15, 'sp4_r_v_b_33')
// (18, 16, 'neigh_op_rgt_2')
// (18, 16, 'sp4_r_v_b_20')
// (18, 17, 'neigh_op_bnr_2')
// (18, 17, 'sp4_r_v_b_9')
// (19, 13, 'sp4_h_r_2')
// (19, 13, 'sp4_v_t_44')
// (19, 14, 'sp4_v_b_44')
// (19, 15, 'neigh_op_top_2')
// (19, 15, 'sp4_v_b_33')
// (19, 16, 'lutff_2/out')
// (19, 16, 'sp4_v_b_20')
// (19, 17, 'neigh_op_bot_2')
// (19, 17, 'sp4_v_b_9')
// (20, 13, 'sp4_h_r_15')
// (20, 15, 'neigh_op_tnl_2')
// (20, 16, 'neigh_op_lft_2')
// (20, 17, 'neigh_op_bnl_2')
// (21, 13, 'local_g2_2')
// (21, 13, 'lutff_1/in_1')
// (21, 13, 'sp4_h_r_26')
// (22, 13, 'sp4_h_r_39')
// (23, 13, 'sp4_h_l_39')

reg n1332 = 0;
// (18, 15, 'local_g2_0')
// (18, 15, 'lutff_4/in_0')
// (18, 15, 'neigh_op_tnr_0')
// (18, 16, 'neigh_op_rgt_0')
// (18, 17, 'neigh_op_bnr_0')
// (19, 15, 'neigh_op_top_0')
// (19, 16, 'lutff_0/out')
// (19, 17, 'neigh_op_bot_0')
// (20, 15, 'neigh_op_tnl_0')
// (20, 16, 'neigh_op_lft_0')
// (20, 17, 'neigh_op_bnl_0')

wire n1333;
// (18, 15, 'lutff_2/lout')
// (18, 15, 'lutff_3/in_2')

wire n1334;
// (18, 15, 'lutff_4/lout')
// (18, 15, 'lutff_5/in_2')

wire n1335;
// (18, 15, 'lutff_5/lout')
// (18, 15, 'lutff_6/in_2')

reg n1336 = 0;
// (18, 15, 'neigh_op_tnr_3')
// (18, 16, 'neigh_op_rgt_3')
// (18, 16, 'sp4_h_r_11')
// (18, 17, 'neigh_op_bnr_3')
// (19, 15, 'neigh_op_top_3')
// (19, 16, 'lutff_3/out')
// (19, 16, 'sp4_h_r_22')
// (19, 17, 'neigh_op_bot_3')
// (20, 15, 'neigh_op_tnl_3')
// (20, 16, 'neigh_op_lft_3')
// (20, 16, 'sp4_h_r_35')
// (20, 17, 'neigh_op_bnl_3')
// (21, 16, 'local_g2_6')
// (21, 16, 'lutff_5/in_1')
// (21, 16, 'sp4_h_r_46')
// (22, 16, 'sp4_h_l_46')

reg n1337 = 0;
// (18, 15, 'neigh_op_tnr_4')
// (18, 16, 'neigh_op_rgt_4')
// (18, 17, 'neigh_op_bnr_4')
// (19, 15, 'neigh_op_top_4')
// (19, 16, 'lutff_4/out')
// (19, 16, 'sp12_h_r_0')
// (19, 17, 'neigh_op_bot_4')
// (20, 15, 'neigh_op_tnl_4')
// (20, 16, 'neigh_op_lft_4')
// (20, 16, 'sp12_h_r_3')
// (20, 17, 'neigh_op_bnl_4')
// (21, 16, 'sp12_h_r_4')
// (22, 16, 'local_g1_7')
// (22, 16, 'lutff_3/in_1')
// (22, 16, 'sp12_h_r_7')
// (23, 16, 'sp12_h_r_8')
// (24, 16, 'sp12_h_r_11')
// (25, 16, 'sp12_h_r_12')
// (26, 16, 'sp12_h_r_15')
// (27, 16, 'sp12_h_r_16')
// (28, 16, 'sp12_h_r_19')
// (29, 16, 'sp12_h_r_20')
// (30, 16, 'sp12_h_r_23')
// (31, 16, 'sp12_h_l_23')

reg n1338 = 0;
// (18, 15, 'neigh_op_tnr_5')
// (18, 16, 'neigh_op_rgt_5')
// (18, 16, 'sp4_r_v_b_42')
// (18, 17, 'neigh_op_bnr_5')
// (18, 17, 'sp4_r_v_b_31')
// (18, 18, 'sp4_r_v_b_18')
// (18, 19, 'sp4_r_v_b_7')
// (19, 15, 'neigh_op_top_5')
// (19, 15, 'sp4_v_t_42')
// (19, 16, 'lutff_5/out')
// (19, 16, 'sp4_v_b_42')
// (19, 17, 'neigh_op_bot_5')
// (19, 17, 'sp4_v_b_31')
// (19, 18, 'local_g0_2')
// (19, 18, 'lutff_7/in_1')
// (19, 18, 'sp4_v_b_18')
// (19, 19, 'sp4_v_b_7')
// (20, 15, 'neigh_op_tnl_5')
// (20, 16, 'neigh_op_lft_5')
// (20, 17, 'neigh_op_bnl_5')

reg n1339 = 0;
// (18, 15, 'neigh_op_tnr_6')
// (18, 15, 'sp4_r_v_b_41')
// (18, 16, 'neigh_op_rgt_6')
// (18, 16, 'sp4_r_v_b_28')
// (18, 17, 'neigh_op_bnr_6')
// (18, 17, 'sp4_r_v_b_17')
// (18, 18, 'sp4_r_v_b_4')
// (19, 14, 'local_g0_4')
// (19, 14, 'lutff_7/in_1')
// (19, 14, 'sp4_h_r_4')
// (19, 14, 'sp4_v_t_41')
// (19, 15, 'neigh_op_top_6')
// (19, 15, 'sp4_v_b_41')
// (19, 16, 'lutff_6/out')
// (19, 16, 'sp4_v_b_28')
// (19, 17, 'neigh_op_bot_6')
// (19, 17, 'sp4_v_b_17')
// (19, 18, 'sp4_v_b_4')
// (20, 14, 'sp4_h_r_17')
// (20, 15, 'neigh_op_tnl_6')
// (20, 16, 'neigh_op_lft_6')
// (20, 17, 'neigh_op_bnl_6')
// (21, 14, 'sp4_h_r_28')
// (22, 14, 'sp4_h_r_41')
// (23, 14, 'sp4_h_l_41')

reg n1340 = 0;
// (18, 15, 'sp12_h_r_1')
// (19, 15, 'local_g0_2')
// (19, 15, 'lutff_3/in_3')
// (19, 15, 'sp12_h_r_2')
// (20, 15, 'sp12_h_r_5')
// (21, 15, 'sp12_h_r_6')
// (22, 14, 'neigh_op_tnr_1')
// (22, 15, 'neigh_op_rgt_1')
// (22, 15, 'sp12_h_r_9')
// (22, 16, 'neigh_op_bnr_1')
// (23, 14, 'neigh_op_top_1')
// (23, 15, 'lutff_1/out')
// (23, 15, 'sp12_h_r_10')
// (23, 16, 'neigh_op_bot_1')
// (24, 14, 'neigh_op_tnl_1')
// (24, 15, 'neigh_op_lft_1')
// (24, 15, 'sp12_h_r_13')
// (24, 16, 'neigh_op_bnl_1')
// (25, 15, 'sp12_h_r_14')
// (26, 15, 'sp12_h_r_17')
// (27, 15, 'sp12_h_r_18')
// (28, 15, 'sp12_h_r_21')
// (29, 15, 'sp12_h_r_22')
// (30, 15, 'sp12_h_l_22')

reg n1341 = 0;
// (18, 15, 'sp4_r_v_b_46')
// (18, 16, 'sp4_r_v_b_35')
// (18, 17, 'sp4_r_v_b_22')
// (18, 18, 'sp4_r_v_b_11')
// (19, 14, 'sp4_h_r_5')
// (19, 14, 'sp4_v_t_46')
// (19, 15, 'sp4_v_b_46')
// (19, 16, 'sp4_v_b_35')
// (19, 17, 'sp4_v_b_22')
// (19, 18, 'local_g1_3')
// (19, 18, 'lutff_1/in_3')
// (19, 18, 'sp4_v_b_11')
// (20, 14, 'sp4_h_r_16')
// (21, 13, 'neigh_op_tnr_4')
// (21, 14, 'neigh_op_rgt_4')
// (21, 14, 'sp4_h_r_29')
// (21, 15, 'neigh_op_bnr_4')
// (22, 13, 'neigh_op_top_4')
// (22, 14, 'lutff_4/out')
// (22, 14, 'sp4_h_r_40')
// (22, 15, 'neigh_op_bot_4')
// (23, 13, 'neigh_op_tnl_4')
// (23, 14, 'neigh_op_lft_4')
// (23, 14, 'sp4_h_l_40')
// (23, 15, 'neigh_op_bnl_4')

wire n1342;
// (18, 16, 'lutff_0/cout')
// (18, 16, 'lutff_1/in_3')

wire n1343;
// (18, 16, 'lutff_1/cout')
// (18, 16, 'lutff_2/in_3')

wire n1344;
// (18, 16, 'lutff_2/cout')
// (18, 16, 'lutff_3/in_3')

wire n1345;
// (18, 16, 'lutff_3/cout')
// (18, 16, 'lutff_4/in_3')

wire n1346;
// (18, 16, 'neigh_op_tnr_3')
// (18, 17, 'neigh_op_rgt_3')
// (18, 18, 'neigh_op_bnr_3')
// (19, 16, 'neigh_op_top_3')
// (19, 17, 'local_g0_3')
// (19, 17, 'lutff_0/in_3')
// (19, 17, 'lutff_3/out')
// (19, 18, 'neigh_op_bot_3')
// (20, 16, 'neigh_op_tnl_3')
// (20, 17, 'neigh_op_lft_3')
// (20, 18, 'neigh_op_bnl_3')

wire n1347;
// (18, 16, 'neigh_op_tnr_6')
// (18, 17, 'neigh_op_rgt_6')
// (18, 18, 'neigh_op_bnr_6')
// (19, 16, 'neigh_op_top_6')
// (19, 17, 'local_g2_6')
// (19, 17, 'lutff_1/in_3')
// (19, 17, 'lutff_6/out')
// (19, 18, 'neigh_op_bot_6')
// (20, 16, 'neigh_op_tnl_6')
// (20, 17, 'neigh_op_lft_6')
// (20, 18, 'neigh_op_bnl_6')

wire n1348;
// (18, 16, 'sp4_r_v_b_36')
// (18, 17, 'sp4_r_v_b_25')
// (18, 18, 'sp4_r_v_b_12')
// (18, 19, 'sp4_r_v_b_1')
// (19, 15, 'sp4_v_t_36')
// (19, 16, 'sp4_v_b_36')
// (19, 17, 'local_g3_1')
// (19, 17, 'lutff_5/in_3')
// (19, 17, 'sp4_v_b_25')
// (19, 18, 'sp4_v_b_12')
// (19, 19, 'sp4_h_r_1')
// (19, 19, 'sp4_v_b_1')
// (20, 19, 'sp4_h_r_12')
// (21, 18, 'neigh_op_tnr_2')
// (21, 19, 'neigh_op_rgt_2')
// (21, 19, 'sp4_h_r_25')
// (21, 20, 'neigh_op_bnr_2')
// (22, 18, 'neigh_op_top_2')
// (22, 19, 'lutff_2/out')
// (22, 19, 'sp4_h_r_36')
// (22, 20, 'neigh_op_bot_2')
// (23, 18, 'neigh_op_tnl_2')
// (23, 19, 'neigh_op_lft_2')
// (23, 19, 'sp4_h_l_36')
// (23, 20, 'neigh_op_bnl_2')

wire n1349;
// (18, 16, 'sp4_r_v_b_43')
// (18, 17, 'sp4_r_v_b_30')
// (18, 18, 'sp4_r_v_b_19')
// (18, 19, 'sp4_r_v_b_6')
// (18, 20, 'sp4_r_v_b_44')
// (18, 21, 'sp4_r_v_b_33')
// (18, 22, 'sp4_r_v_b_20')
// (18, 23, 'sp4_r_v_b_9')
// (19, 15, 'sp4_h_r_6')
// (19, 15, 'sp4_v_t_43')
// (19, 16, 'sp4_v_b_43')
// (19, 17, 'sp4_v_b_30')
// (19, 18, 'sp4_v_b_19')
// (19, 19, 'sp4_v_b_6')
// (19, 19, 'sp4_v_t_44')
// (19, 20, 'sp4_v_b_44')
// (19, 21, 'local_g3_1')
// (19, 21, 'lutff_5/in_1')
// (19, 21, 'sp4_v_b_33')
// (19, 22, 'sp4_v_b_20')
// (19, 23, 'sp4_v_b_9')
// (20, 15, 'sp4_h_r_19')
// (21, 15, 'sp4_h_r_30')
// (22, 15, 'sp12_h_r_0')
// (22, 15, 'sp4_h_r_43')
// (23, 15, 'sp12_h_r_3')
// (23, 15, 'sp4_h_l_43')
// (23, 15, 'sp4_h_r_3')
// (24, 15, 'sp12_h_r_4')
// (24, 15, 'sp4_h_r_14')
// (25, 15, 'sp12_h_r_7')
// (25, 15, 'sp4_h_r_27')
// (26, 15, 'sp12_h_r_8')
// (26, 15, 'sp4_h_r_38')
// (27, 15, 'sp12_h_r_11')
// (27, 15, 'sp4_h_l_38')
// (28, 15, 'sp12_h_r_12')
// (29, 15, 'sp12_h_r_15')
// (30, 15, 'sp12_h_r_16')
// (31, 15, 'sp12_h_r_19')
// (32, 14, 'neigh_op_tnr_2')
// (32, 14, 'neigh_op_tnr_6')
// (32, 15, 'neigh_op_rgt_2')
// (32, 15, 'neigh_op_rgt_6')
// (32, 15, 'sp12_h_r_20')
// (32, 16, 'neigh_op_bnr_2')
// (32, 16, 'neigh_op_bnr_6')
// (33, 15, 'io_1/D_IN_0')
// (33, 15, 'span12_horz_20')

wire n1350;
// (18, 16, 'sp4_r_v_b_44')
// (18, 17, 'local_g2_1')
// (18, 17, 'lutff_6/in_3')
// (18, 17, 'sp4_r_v_b_33')
// (18, 18, 'sp4_r_v_b_20')
// (18, 19, 'sp4_r_v_b_9')
// (19, 15, 'sp4_v_t_44')
// (19, 16, 'sp4_v_b_44')
// (19, 17, 'sp4_v_b_33')
// (19, 18, 'sp4_v_b_20')
// (19, 19, 'sp4_h_r_9')
// (19, 19, 'sp4_v_b_9')
// (20, 19, 'sp4_h_r_20')
// (21, 18, 'neigh_op_tnr_6')
// (21, 19, 'neigh_op_rgt_6')
// (21, 19, 'sp4_h_r_33')
// (21, 20, 'neigh_op_bnr_6')
// (22, 18, 'neigh_op_top_6')
// (22, 19, 'lutff_6/out')
// (22, 19, 'sp4_h_r_44')
// (22, 20, 'neigh_op_bot_6')
// (23, 18, 'neigh_op_tnl_6')
// (23, 19, 'neigh_op_lft_6')
// (23, 19, 'sp4_h_l_44')
// (23, 20, 'neigh_op_bnl_6')

reg n1351 = 0;
// (18, 17, 'local_g0_4')
// (18, 17, 'lutff_7/in_3')
// (18, 17, 'sp4_h_r_4')
// (19, 17, 'sp4_h_r_17')
// (20, 17, 'sp4_h_r_28')
// (21, 17, 'sp4_h_r_41')
// (21, 18, 'sp4_r_v_b_41')
// (21, 19, 'sp4_r_v_b_28')
// (21, 20, 'sp4_r_v_b_17')
// (21, 21, 'sp4_r_v_b_4')
// (21, 22, 'neigh_op_tnr_0')
// (21, 22, 'sp4_r_v_b_45')
// (21, 23, 'neigh_op_rgt_0')
// (21, 23, 'sp4_r_v_b_32')
// (21, 24, 'neigh_op_bnr_0')
// (21, 24, 'sp4_r_v_b_21')
// (21, 25, 'sp4_r_v_b_8')
// (22, 17, 'sp4_h_l_41')
// (22, 17, 'sp4_v_t_41')
// (22, 18, 'sp4_v_b_41')
// (22, 19, 'sp4_v_b_28')
// (22, 20, 'sp4_v_b_17')
// (22, 21, 'sp4_v_b_4')
// (22, 21, 'sp4_v_t_45')
// (22, 22, 'neigh_op_top_0')
// (22, 22, 'sp4_v_b_45')
// (22, 23, 'lutff_0/out')
// (22, 23, 'sp4_v_b_32')
// (22, 24, 'neigh_op_bot_0')
// (22, 24, 'sp4_v_b_21')
// (22, 25, 'sp4_v_b_8')
// (23, 22, 'neigh_op_tnl_0')
// (23, 23, 'neigh_op_lft_0')
// (23, 24, 'neigh_op_bnl_0')

wire n1352;
// (18, 17, 'lutff_1/lout')
// (18, 17, 'lutff_2/in_2')

wire n1353;
// (18, 17, 'lutff_4/lout')
// (18, 17, 'lutff_5/in_2')

wire n1354;
// (18, 17, 'lutff_5/lout')
// (18, 17, 'lutff_6/in_2')

reg n1355 = 0;
// (18, 17, 'neigh_op_tnr_0')
// (18, 18, 'neigh_op_rgt_0')
// (18, 19, 'neigh_op_bnr_0')
// (19, 17, 'neigh_op_top_0')
// (19, 18, 'local_g1_0')
// (19, 18, 'lutff_0/out')
// (19, 18, 'lutff_2/in_3')
// (19, 19, 'neigh_op_bot_0')
// (20, 17, 'neigh_op_tnl_0')
// (20, 18, 'neigh_op_lft_0')
// (20, 19, 'neigh_op_bnl_0')

wire n1356;
// (18, 17, 'neigh_op_tnr_2')
// (18, 18, 'neigh_op_rgt_2')
// (18, 19, 'neigh_op_bnr_2')
// (19, 17, 'neigh_op_top_2')
// (19, 18, 'lutff_2/out')
// (19, 18, 'sp4_h_r_4')
// (19, 19, 'neigh_op_bot_2')
// (20, 17, 'neigh_op_tnl_2')
// (20, 18, 'neigh_op_lft_2')
// (20, 18, 'sp4_h_r_17')
// (20, 19, 'neigh_op_bnl_2')
// (21, 18, 'sp4_h_r_28')
// (22, 18, 'local_g3_1')
// (22, 18, 'lutff_3/in_1')
// (22, 18, 'sp4_h_r_41')
// (23, 18, 'sp4_h_l_41')

wire n1357;
// (18, 17, 'neigh_op_tnr_5')
// (18, 18, 'neigh_op_rgt_5')
// (18, 19, 'neigh_op_bnr_5')
// (19, 17, 'local_g1_5')
// (19, 17, 'lutff_1/in_1')
// (19, 17, 'neigh_op_top_5')
// (19, 18, 'lutff_5/out')
// (19, 19, 'neigh_op_bot_5')
// (20, 17, 'neigh_op_tnl_5')
// (20, 18, 'neigh_op_lft_5')
// (20, 19, 'neigh_op_bnl_5')

wire n1358;
// (18, 17, 'neigh_op_tnr_6')
// (18, 18, 'neigh_op_rgt_6')
// (18, 19, 'neigh_op_bnr_6')
// (19, 17, 'neigh_op_top_6')
// (19, 18, 'local_g2_6')
// (19, 18, 'lutff_5/in_3')
// (19, 18, 'lutff_6/out')
// (19, 19, 'neigh_op_bot_6')
// (20, 17, 'neigh_op_tnl_6')
// (20, 18, 'neigh_op_lft_6')
// (20, 19, 'neigh_op_bnl_6')

wire n1359;
// (18, 17, 'neigh_op_tnr_7')
// (18, 18, 'neigh_op_rgt_7')
// (18, 19, 'neigh_op_bnr_7')
// (19, 17, 'neigh_op_top_7')
// (19, 18, 'local_g2_7')
// (19, 18, 'lutff_6/in_3')
// (19, 18, 'lutff_7/out')
// (19, 19, 'neigh_op_bot_7')
// (20, 17, 'neigh_op_tnl_7')
// (20, 18, 'neigh_op_lft_7')
// (20, 19, 'neigh_op_bnl_7')

reg n1360 = 0;
// (18, 17, 'sp12_h_r_0')
// (19, 17, 'sp12_h_r_3')
// (20, 17, 'local_g1_4')
// (20, 17, 'lutff_4/in_1')
// (20, 17, 'sp12_h_r_4')
// (21, 17, 'sp12_h_r_7')
// (22, 17, 'sp12_h_r_8')
// (23, 16, 'neigh_op_tnr_2')
// (23, 17, 'neigh_op_rgt_2')
// (23, 17, 'sp12_h_r_11')
// (23, 18, 'neigh_op_bnr_2')
// (24, 16, 'neigh_op_top_2')
// (24, 17, 'lutff_2/out')
// (24, 17, 'sp12_h_r_12')
// (24, 18, 'neigh_op_bot_2')
// (25, 16, 'neigh_op_tnl_2')
// (25, 17, 'neigh_op_lft_2')
// (25, 17, 'sp12_h_r_15')
// (25, 18, 'neigh_op_bnl_2')
// (26, 17, 'sp12_h_r_16')
// (27, 17, 'sp12_h_r_19')
// (28, 17, 'sp12_h_r_20')
// (29, 17, 'sp12_h_r_23')
// (30, 17, 'sp12_h_l_23')

reg n1361 = 0;
// (18, 18, 'local_g1_0')
// (18, 18, 'lutff_4/in_3')
// (18, 18, 'sp4_h_r_0')
// (19, 18, 'sp4_h_r_13')
// (20, 18, 'sp4_h_r_24')
// (21, 18, 'sp4_h_r_37')
// (21, 19, 'sp4_r_v_b_37')
// (21, 20, 'sp4_r_v_b_24')
// (21, 21, 'sp4_r_v_b_13')
// (21, 22, 'neigh_op_tnr_6')
// (21, 22, 'sp4_r_v_b_0')
// (21, 23, 'neigh_op_rgt_6')
// (21, 23, 'sp4_r_v_b_44')
// (21, 24, 'neigh_op_bnr_6')
// (21, 24, 'sp4_r_v_b_33')
// (21, 25, 'sp4_r_v_b_20')
// (21, 26, 'sp4_r_v_b_9')
// (22, 18, 'sp4_h_l_37')
// (22, 18, 'sp4_v_t_37')
// (22, 19, 'sp4_v_b_37')
// (22, 20, 'sp4_v_b_24')
// (22, 21, 'sp4_v_b_13')
// (22, 22, 'neigh_op_top_6')
// (22, 22, 'sp4_v_b_0')
// (22, 22, 'sp4_v_t_44')
// (22, 23, 'lutff_6/out')
// (22, 23, 'sp4_v_b_44')
// (22, 24, 'neigh_op_bot_6')
// (22, 24, 'sp4_v_b_33')
// (22, 25, 'sp4_v_b_20')
// (22, 26, 'sp4_v_b_9')
// (23, 22, 'neigh_op_tnl_6')
// (23, 23, 'neigh_op_lft_6')
// (23, 24, 'neigh_op_bnl_6')

reg n1362 = 0;
// (18, 18, 'local_g2_5')
// (18, 18, 'lutff_1/in_0')
// (18, 18, 'sp4_r_v_b_37')
// (18, 19, 'sp4_r_v_b_24')
// (18, 20, 'sp4_r_v_b_13')
// (18, 21, 'sp4_r_v_b_0')
// (19, 17, 'sp4_v_t_37')
// (19, 18, 'sp4_v_b_37')
// (19, 19, 'sp4_v_b_24')
// (19, 20, 'sp4_v_b_13')
// (19, 21, 'sp4_h_r_7')
// (19, 21, 'sp4_v_b_0')
// (20, 21, 'sp4_h_r_18')
// (21, 20, 'neigh_op_tnr_5')
// (21, 21, 'neigh_op_rgt_5')
// (21, 21, 'sp4_h_r_31')
// (21, 22, 'neigh_op_bnr_5')
// (22, 20, 'neigh_op_top_5')
// (22, 21, 'lutff_5/out')
// (22, 21, 'sp4_h_r_42')
// (22, 22, 'neigh_op_bot_5')
// (23, 20, 'neigh_op_tnl_5')
// (23, 21, 'neigh_op_lft_5')
// (23, 21, 'sp4_h_l_42')
// (23, 22, 'neigh_op_bnl_5')

wire n1363;
// (18, 18, 'lutff_1/lout')
// (18, 18, 'lutff_2/in_2')

wire n1364;
// (18, 18, 'lutff_5/lout')
// (18, 18, 'lutff_6/in_2')

wire n1365;
// (18, 18, 'lutff_6/lout')
// (18, 18, 'lutff_7/in_2')

reg n1366 = 0;
// (18, 18, 'neigh_op_tnr_1')
// (18, 19, 'neigh_op_rgt_1')
// (18, 19, 'sp4_h_r_7')
// (18, 20, 'neigh_op_bnr_1')
// (19, 18, 'neigh_op_top_1')
// (19, 19, 'lutff_1/out')
// (19, 19, 'sp4_h_r_18')
// (19, 20, 'neigh_op_bot_1')
// (20, 18, 'neigh_op_tnl_1')
// (20, 19, 'neigh_op_lft_1')
// (20, 19, 'sp4_h_r_31')
// (20, 20, 'neigh_op_bnl_1')
// (21, 16, 'sp4_r_v_b_36')
// (21, 17, 'sp4_r_v_b_25')
// (21, 18, 'local_g2_4')
// (21, 18, 'lutff_1/in_3')
// (21, 18, 'sp4_r_v_b_12')
// (21, 19, 'sp4_h_r_42')
// (21, 19, 'sp4_r_v_b_1')
// (22, 15, 'sp4_v_t_36')
// (22, 16, 'sp4_v_b_36')
// (22, 17, 'sp4_v_b_25')
// (22, 18, 'sp4_v_b_12')
// (22, 19, 'sp4_h_l_42')
// (22, 19, 'sp4_v_b_1')

reg n1367 = 0;
// (18, 18, 'neigh_op_tnr_2')
// (18, 19, 'neigh_op_rgt_2')
// (18, 20, 'neigh_op_bnr_2')
// (19, 18, 'neigh_op_top_2')
// (19, 19, 'lutff_2/out')
// (19, 19, 'sp4_r_v_b_37')
// (19, 20, 'neigh_op_bot_2')
// (19, 20, 'sp4_r_v_b_24')
// (19, 21, 'sp4_r_v_b_13')
// (19, 22, 'sp4_r_v_b_0')
// (20, 18, 'neigh_op_tnl_2')
// (20, 18, 'sp4_h_r_5')
// (20, 18, 'sp4_v_t_37')
// (20, 19, 'neigh_op_lft_2')
// (20, 19, 'sp4_v_b_37')
// (20, 20, 'neigh_op_bnl_2')
// (20, 20, 'sp4_v_b_24')
// (20, 21, 'sp4_v_b_13')
// (20, 22, 'sp4_v_b_0')
// (21, 18, 'local_g1_0')
// (21, 18, 'lutff_4/in_3')
// (21, 18, 'sp4_h_r_16')
// (22, 18, 'sp4_h_r_29')
// (23, 18, 'sp4_h_r_40')
// (24, 18, 'sp4_h_l_40')

reg n1368 = 0;
// (18, 18, 'neigh_op_tnr_3')
// (18, 19, 'neigh_op_rgt_3')
// (18, 19, 'sp4_r_v_b_38')
// (18, 20, 'neigh_op_bnr_3')
// (18, 20, 'sp4_r_v_b_27')
// (18, 21, 'sp4_r_v_b_14')
// (18, 22, 'sp4_r_v_b_3')
// (19, 18, 'neigh_op_top_3')
// (19, 18, 'sp4_h_r_3')
// (19, 18, 'sp4_v_t_38')
// (19, 19, 'lutff_3/out')
// (19, 19, 'sp4_v_b_38')
// (19, 20, 'neigh_op_bot_3')
// (19, 20, 'sp4_v_b_27')
// (19, 21, 'sp4_v_b_14')
// (19, 22, 'sp4_v_b_3')
// (20, 18, 'neigh_op_tnl_3')
// (20, 18, 'sp4_h_r_14')
// (20, 19, 'neigh_op_lft_3')
// (20, 20, 'neigh_op_bnl_3')
// (21, 18, 'local_g3_3')
// (21, 18, 'lutff_7/in_3')
// (21, 18, 'sp4_h_r_27')
// (22, 18, 'sp4_h_r_38')
// (23, 18, 'sp4_h_l_38')

wire n1369;
// (18, 18, 'sp4_h_r_1')
// (18, 18, 'sp4_h_r_10')
// (19, 18, 'sp4_h_r_12')
// (19, 18, 'sp4_h_r_23')
// (20, 18, 'local_g2_2')
// (20, 18, 'lutff_global/cen')
// (20, 18, 'sp4_h_r_25')
// (20, 18, 'sp4_h_r_34')
// (21, 14, 'neigh_op_tnr_2')
// (21, 15, 'neigh_op_rgt_2')
// (21, 15, 'sp4_r_v_b_36')
// (21, 16, 'neigh_op_bnr_2')
// (21, 16, 'sp4_r_v_b_25')
// (21, 17, 'sp4_r_v_b_12')
// (21, 18, 'sp4_h_r_36')
// (21, 18, 'sp4_h_r_47')
// (21, 18, 'sp4_r_v_b_1')
// (21, 19, 'sp4_r_v_b_41')
// (21, 19, 'sp4_r_v_b_43')
// (21, 20, 'sp4_r_v_b_28')
// (21, 20, 'sp4_r_v_b_30')
// (21, 21, 'sp4_r_v_b_17')
// (21, 21, 'sp4_r_v_b_19')
// (21, 22, 'sp4_r_v_b_4')
// (21, 22, 'sp4_r_v_b_6')
// (22, 13, 'sp12_v_t_23')
// (22, 14, 'neigh_op_top_2')
// (22, 14, 'sp12_v_b_23')
// (22, 14, 'sp4_v_t_36')
// (22, 15, 'lutff_2/out')
// (22, 15, 'sp12_v_b_20')
// (22, 15, 'sp4_v_b_36')
// (22, 16, 'neigh_op_bot_2')
// (22, 16, 'sp12_v_b_19')
// (22, 16, 'sp4_v_b_25')
// (22, 17, 'sp12_v_b_16')
// (22, 17, 'sp4_v_b_12')
// (22, 18, 'sp12_v_b_15')
// (22, 18, 'sp4_h_l_36')
// (22, 18, 'sp4_h_l_47')
// (22, 18, 'sp4_v_b_1')
// (22, 18, 'sp4_v_t_41')
// (22, 18, 'sp4_v_t_43')
// (22, 19, 'local_g3_3')
// (22, 19, 'lutff_global/cen')
// (22, 19, 'sp12_v_b_12')
// (22, 19, 'sp4_v_b_41')
// (22, 19, 'sp4_v_b_43')
// (22, 20, 'sp12_v_b_11')
// (22, 20, 'sp4_v_b_28')
// (22, 20, 'sp4_v_b_30')
// (22, 21, 'sp12_v_b_8')
// (22, 21, 'sp4_v_b_17')
// (22, 21, 'sp4_v_b_19')
// (22, 22, 'sp12_v_b_7')
// (22, 22, 'sp4_v_b_4')
// (22, 22, 'sp4_v_b_6')
// (22, 23, 'sp12_v_b_4')
// (22, 24, 'local_g3_3')
// (22, 24, 'lutff_global/cen')
// (22, 24, 'sp12_v_b_3')
// (22, 25, 'sp12_v_b_0')
// (23, 14, 'neigh_op_tnl_2')
// (23, 15, 'neigh_op_lft_2')
// (23, 16, 'neigh_op_bnl_2')

reg n1370 = 0;
// (18, 18, 'sp4_h_r_8')
// (19, 18, 'local_g1_5')
// (19, 18, 'lutff_3/in_3')
// (19, 18, 'sp4_h_r_21')
// (20, 18, 'sp4_h_r_32')
// (21, 15, 'sp4_r_v_b_45')
// (21, 16, 'sp4_r_v_b_32')
// (21, 17, 'sp4_r_v_b_21')
// (21, 18, 'sp4_h_r_45')
// (21, 18, 'sp4_r_v_b_8')
// (22, 14, 'sp4_h_r_2')
// (22, 14, 'sp4_v_t_45')
// (22, 15, 'sp4_v_b_45')
// (22, 16, 'sp4_v_b_32')
// (22, 17, 'sp4_v_b_21')
// (22, 18, 'sp4_h_l_45')
// (22, 18, 'sp4_v_b_8')
// (23, 13, 'neigh_op_tnr_5')
// (23, 14, 'neigh_op_rgt_5')
// (23, 14, 'sp4_h_r_15')
// (23, 15, 'neigh_op_bnr_5')
// (24, 13, 'neigh_op_top_5')
// (24, 14, 'lutff_5/out')
// (24, 14, 'sp4_h_r_26')
// (24, 15, 'neigh_op_bot_5')
// (25, 13, 'neigh_op_tnl_5')
// (25, 14, 'neigh_op_lft_5')
// (25, 14, 'sp4_h_r_39')
// (25, 15, 'neigh_op_bnl_5')
// (26, 14, 'sp4_h_l_39')

reg n1371 = 0;
// (18, 19, 'local_g1_0')
// (18, 19, 'lutff_2/in_3')
// (18, 19, 'sp4_h_r_8')
// (19, 18, 'neigh_op_tnr_0')
// (19, 19, 'neigh_op_rgt_0')
// (19, 19, 'sp4_h_r_21')
// (19, 20, 'neigh_op_bnr_0')
// (20, 18, 'neigh_op_top_0')
// (20, 19, 'lutff_0/out')
// (20, 19, 'sp4_h_r_32')
// (20, 20, 'neigh_op_bot_0')
// (21, 18, 'neigh_op_tnl_0')
// (21, 19, 'neigh_op_lft_0')
// (21, 19, 'sp4_h_r_45')
// (21, 20, 'neigh_op_bnl_0')
// (22, 19, 'sp4_h_l_45')

reg n1372 = 0;
// (18, 19, 'local_g1_2')
// (18, 19, 'lutff_0/in_1')
// (18, 19, 'sp4_h_r_10')
// (19, 19, 'sp4_h_r_23')
// (20, 19, 'sp4_h_r_34')
// (21, 19, 'sp4_h_r_47')
// (21, 20, 'neigh_op_tnr_6')
// (21, 20, 'sp4_r_v_b_41')
// (21, 21, 'neigh_op_rgt_6')
// (21, 21, 'sp4_r_v_b_28')
// (21, 22, 'neigh_op_bnr_6')
// (21, 22, 'sp4_r_v_b_17')
// (21, 23, 'sp4_r_v_b_4')
// (22, 19, 'sp4_h_l_47')
// (22, 19, 'sp4_v_t_41')
// (22, 20, 'neigh_op_top_6')
// (22, 20, 'sp4_v_b_41')
// (22, 21, 'lutff_6/out')
// (22, 21, 'sp4_v_b_28')
// (22, 22, 'neigh_op_bot_6')
// (22, 22, 'sp4_v_b_17')
// (22, 23, 'sp4_v_b_4')
// (23, 20, 'neigh_op_tnl_6')
// (23, 21, 'neigh_op_lft_6')
// (23, 22, 'neigh_op_bnl_6')

reg n1373 = 0;
// (18, 19, 'local_g1_4')
// (18, 19, 'lutff_4/in_3')
// (18, 19, 'sp4_h_r_4')
// (19, 18, 'neigh_op_tnr_6')
// (19, 19, 'neigh_op_rgt_6')
// (19, 19, 'sp4_h_r_17')
// (19, 20, 'neigh_op_bnr_6')
// (20, 18, 'neigh_op_top_6')
// (20, 19, 'lutff_6/out')
// (20, 19, 'sp4_h_r_28')
// (20, 20, 'neigh_op_bot_6')
// (21, 18, 'neigh_op_tnl_6')
// (21, 19, 'neigh_op_lft_6')
// (21, 19, 'sp4_h_r_41')
// (21, 20, 'neigh_op_bnl_6')
// (22, 19, 'sp4_h_l_41')

reg n1374 = 0;
// (18, 19, 'local_g2_4')
// (18, 19, 'lutff_5/in_3')
// (18, 19, 'sp4_r_v_b_36')
// (18, 20, 'sp4_r_v_b_25')
// (18, 21, 'sp4_r_v_b_12')
// (18, 22, 'sp4_r_v_b_1')
// (18, 23, 'sp4_r_v_b_40')
// (18, 24, 'neigh_op_tnr_0')
// (18, 24, 'sp4_r_v_b_29')
// (18, 25, 'neigh_op_rgt_0')
// (18, 25, 'sp4_r_v_b_16')
// (18, 26, 'neigh_op_bnr_0')
// (18, 26, 'sp4_r_v_b_5')
// (19, 18, 'sp4_v_t_36')
// (19, 19, 'sp4_v_b_36')
// (19, 20, 'sp4_v_b_25')
// (19, 21, 'sp4_v_b_12')
// (19, 22, 'sp4_v_b_1')
// (19, 22, 'sp4_v_t_40')
// (19, 23, 'sp4_v_b_40')
// (19, 24, 'neigh_op_top_0')
// (19, 24, 'sp4_v_b_29')
// (19, 25, 'lutff_0/out')
// (19, 25, 'sp4_v_b_16')
// (19, 26, 'neigh_op_bot_0')
// (19, 26, 'sp4_v_b_5')
// (20, 24, 'neigh_op_tnl_0')
// (20, 25, 'neigh_op_lft_0')
// (20, 26, 'neigh_op_bnl_0')

reg n1375 = 0;
// (18, 19, 'local_g3_2')
// (18, 19, 'lutff_6/in_3')
// (18, 19, 'sp4_r_v_b_42')
// (18, 20, 'sp4_r_v_b_31')
// (18, 21, 'sp4_r_v_b_18')
// (18, 22, 'sp4_r_v_b_7')
// (18, 23, 'sp4_r_v_b_42')
// (18, 24, 'neigh_op_tnr_1')
// (18, 24, 'sp4_r_v_b_31')
// (18, 25, 'neigh_op_rgt_1')
// (18, 25, 'sp4_r_v_b_18')
// (18, 26, 'neigh_op_bnr_1')
// (18, 26, 'sp4_r_v_b_7')
// (19, 18, 'sp4_v_t_42')
// (19, 19, 'sp4_v_b_42')
// (19, 20, 'sp4_v_b_31')
// (19, 21, 'sp4_v_b_18')
// (19, 22, 'sp4_v_b_7')
// (19, 22, 'sp4_v_t_42')
// (19, 23, 'sp4_v_b_42')
// (19, 24, 'neigh_op_top_1')
// (19, 24, 'sp4_v_b_31')
// (19, 25, 'lutff_1/out')
// (19, 25, 'sp4_v_b_18')
// (19, 26, 'neigh_op_bot_1')
// (19, 26, 'sp4_v_b_7')
// (20, 24, 'neigh_op_tnl_1')
// (20, 25, 'neigh_op_lft_1')
// (20, 26, 'neigh_op_bnl_1')

reg n1376 = 0;
// (18, 19, 'neigh_op_tnr_0')
// (18, 20, 'neigh_op_rgt_0')
// (18, 21, 'neigh_op_bnr_0')
// (19, 8, 'sp12_h_r_0')
// (19, 8, 'sp12_v_t_23')
// (19, 9, 'sp12_v_b_23')
// (19, 10, 'sp12_v_b_20')
// (19, 11, 'sp12_v_b_19')
// (19, 12, 'sp12_v_b_16')
// (19, 13, 'sp12_v_b_15')
// (19, 14, 'sp12_v_b_12')
// (19, 15, 'sp12_v_b_11')
// (19, 16, 'sp12_v_b_8')
// (19, 17, 'sp12_v_b_7')
// (19, 18, 'sp12_v_b_4')
// (19, 19, 'neigh_op_top_0')
// (19, 19, 'sp12_v_b_3')
// (19, 20, 'local_g1_0')
// (19, 20, 'lutff_0/in_1')
// (19, 20, 'lutff_0/out')
// (19, 20, 'sp12_v_b_0')
// (19, 21, 'neigh_op_bot_0')
// (20, 8, 'sp12_h_r_3')
// (20, 19, 'neigh_op_tnl_0')
// (20, 20, 'neigh_op_lft_0')
// (20, 21, 'neigh_op_bnl_0')
// (21, 8, 'sp12_h_r_4')
// (22, 8, 'sp12_h_r_7')
// (23, 8, 'sp12_h_r_8')
// (24, 8, 'sp12_h_r_11')
// (25, 8, 'sp12_h_r_12')
// (26, 8, 'sp12_h_r_15')
// (27, 8, 'sp12_h_r_16')
// (28, 8, 'sp12_h_r_19')
// (29, 8, 'sp12_h_r_20')
// (30, 3, 'sp4_r_v_b_39')
// (30, 4, 'sp4_r_v_b_26')
// (30, 5, 'sp4_r_v_b_15')
// (30, 6, 'sp4_r_v_b_2')
// (30, 8, 'sp12_h_r_23')
// (31, 0, 'span12_vert_15')
// (31, 1, 'sp12_v_b_15')
// (31, 2, 'sp12_v_b_12')
// (31, 2, 'sp4_h_r_7')
// (31, 2, 'sp4_v_t_39')
// (31, 3, 'sp12_v_b_11')
// (31, 3, 'sp4_v_b_39')
// (31, 4, 'sp12_v_b_8')
// (31, 4, 'sp4_v_b_26')
// (31, 5, 'sp12_v_b_7')
// (31, 5, 'sp4_v_b_15')
// (31, 6, 'sp12_v_b_4')
// (31, 6, 'sp4_v_b_2')
// (31, 7, 'sp12_v_b_3')
// (31, 8, 'sp12_h_l_23')
// (31, 8, 'sp12_v_b_0')
// (32, 2, 'sp4_h_r_18')
// (33, 2, 'io_1/OUT_ENB')
// (33, 2, 'local_g0_2')
// (33, 2, 'span4_horz_18')

reg n1377 = 0;
// (18, 19, 'neigh_op_tnr_1')
// (18, 20, 'neigh_op_rgt_1')
// (18, 21, 'neigh_op_bnr_1')
// (19, 9, 'sp12_v_t_22')
// (19, 10, 'sp12_v_b_22')
// (19, 11, 'sp12_v_b_21')
// (19, 12, 'sp12_v_b_18')
// (19, 13, 'sp12_v_b_17')
// (19, 14, 'sp12_v_b_14')
// (19, 15, 'sp12_v_b_13')
// (19, 16, 'sp12_v_b_10')
// (19, 17, 'sp12_v_b_9')
// (19, 18, 'sp12_v_b_6')
// (19, 19, 'neigh_op_top_1')
// (19, 19, 'sp12_v_b_5')
// (19, 20, 'local_g2_1')
// (19, 20, 'lutff_1/in_2')
// (19, 20, 'lutff_1/out')
// (19, 20, 'sp12_v_b_2')
// (19, 21, 'neigh_op_bot_1')
// (19, 21, 'sp12_h_r_1')
// (19, 21, 'sp12_v_b_1')
// (20, 19, 'neigh_op_tnl_1')
// (20, 20, 'neigh_op_lft_1')
// (20, 21, 'neigh_op_bnl_1')
// (20, 21, 'sp12_h_r_2')
// (21, 21, 'sp12_h_r_5')
// (22, 21, 'sp12_h_r_6')
// (23, 21, 'sp12_h_r_9')
// (24, 21, 'sp12_h_r_10')
// (25, 21, 'sp12_h_r_13')
// (26, 21, 'sp12_h_r_14')
// (27, 21, 'sp12_h_r_17')
// (28, 21, 'sp12_h_r_18')
// (29, 21, 'sp12_h_r_21')
// (30, 15, 'sp4_r_v_b_40')
// (30, 16, 'sp4_r_v_b_29')
// (30, 17, 'sp4_r_v_b_16')
// (30, 18, 'sp4_r_v_b_5')
// (30, 21, 'sp12_h_r_22')
// (31, 9, 'sp12_v_t_22')
// (31, 10, 'sp12_v_b_22')
// (31, 11, 'sp12_v_b_21')
// (31, 12, 'sp12_v_b_18')
// (31, 13, 'sp12_v_b_17')
// (31, 14, 'sp12_v_b_14')
// (31, 14, 'sp4_h_r_5')
// (31, 14, 'sp4_v_t_40')
// (31, 15, 'sp12_v_b_13')
// (31, 15, 'sp4_v_b_40')
// (31, 16, 'sp12_v_b_10')
// (31, 16, 'sp4_v_b_29')
// (31, 17, 'sp12_v_b_9')
// (31, 17, 'sp4_v_b_16')
// (31, 18, 'sp12_v_b_6')
// (31, 18, 'sp4_v_b_5')
// (31, 19, 'sp12_v_b_5')
// (31, 20, 'sp12_v_b_2')
// (31, 21, 'sp12_h_l_22')
// (31, 21, 'sp12_v_b_1')
// (32, 14, 'sp4_h_r_16')
// (33, 14, 'io_1/OUT_ENB')
// (33, 14, 'local_g0_0')
// (33, 14, 'span4_horz_16')

reg n1378 = 0;
// (18, 19, 'neigh_op_tnr_2')
// (18, 20, 'neigh_op_rgt_2')
// (18, 21, 'neigh_op_bnr_2')
// (19, 18, 'sp12_v_t_23')
// (19, 19, 'neigh_op_top_2')
// (19, 19, 'sp12_v_b_23')
// (19, 20, 'local_g3_2')
// (19, 20, 'lutff_2/in_1')
// (19, 20, 'lutff_2/out')
// (19, 20, 'sp12_v_b_20')
// (19, 21, 'neigh_op_bot_2')
// (19, 21, 'sp12_v_b_19')
// (19, 22, 'sp12_v_b_16')
// (19, 23, 'sp12_v_b_15')
// (19, 24, 'sp12_v_b_12')
// (19, 25, 'sp12_v_b_11')
// (19, 26, 'sp12_v_b_8')
// (19, 27, 'sp12_v_b_7')
// (19, 28, 'sp12_v_b_4')
// (19, 29, 'sp12_v_b_3')
// (19, 30, 'sp12_h_r_0')
// (19, 30, 'sp12_v_b_0')
// (20, 19, 'neigh_op_tnl_2')
// (20, 20, 'neigh_op_lft_2')
// (20, 21, 'neigh_op_bnl_2')
// (20, 30, 'sp12_h_r_3')
// (21, 30, 'sp12_h_r_4')
// (22, 30, 'sp12_h_r_7')
// (23, 30, 'sp12_h_r_8')
// (24, 30, 'sp12_h_r_11')
// (25, 30, 'sp12_h_r_12')
// (26, 30, 'sp12_h_r_15')
// (26, 30, 'sp4_h_r_9')
// (27, 30, 'sp12_h_r_16')
// (27, 30, 'sp4_h_r_20')
// (28, 30, 'sp12_h_r_19')
// (28, 30, 'sp4_h_r_33')
// (29, 30, 'sp12_h_r_20')
// (29, 30, 'sp4_h_r_44')
// (29, 31, 'sp4_r_v_b_39')
// (29, 32, 'sp4_r_v_b_26')
// (30, 30, 'sp12_h_r_23')
// (30, 30, 'sp4_h_l_44')
// (30, 30, 'sp4_v_t_39')
// (30, 31, 'sp4_v_b_39')
// (30, 32, 'sp4_v_b_26')
// (30, 33, 'io_0/OUT_ENB')
// (30, 33, 'local_g0_7')
// (30, 33, 'span4_vert_15')
// (31, 30, 'sp12_h_l_23')

reg n1379 = 0;
// (18, 19, 'neigh_op_tnr_3')
// (18, 20, 'neigh_op_rgt_3')
// (18, 21, 'neigh_op_bnr_3')
// (19, 19, 'neigh_op_top_3')
// (19, 19, 'sp12_v_t_22')
// (19, 20, 'local_g0_3')
// (19, 20, 'lutff_3/in_2')
// (19, 20, 'lutff_3/out')
// (19, 20, 'sp12_v_b_22')
// (19, 21, 'neigh_op_bot_3')
// (19, 21, 'sp12_v_b_21')
// (19, 22, 'sp12_v_b_18')
// (19, 23, 'sp12_v_b_17')
// (19, 24, 'sp12_v_b_14')
// (19, 25, 'sp12_v_b_13')
// (19, 26, 'sp12_v_b_10')
// (19, 27, 'sp12_v_b_9')
// (19, 28, 'sp12_v_b_6')
// (19, 29, 'sp12_v_b_5')
// (19, 30, 'sp12_v_b_2')
// (19, 31, 'sp12_h_r_1')
// (19, 31, 'sp12_v_b_1')
// (20, 19, 'neigh_op_tnl_3')
// (20, 20, 'neigh_op_lft_3')
// (20, 21, 'neigh_op_bnl_3')
// (20, 31, 'sp12_h_r_2')
// (21, 31, 'sp12_h_r_5')
// (22, 31, 'sp12_h_r_6')
// (23, 31, 'sp12_h_r_9')
// (24, 31, 'sp12_h_r_10')
// (25, 31, 'sp12_h_r_13')
// (26, 31, 'sp12_h_r_14')
// (27, 31, 'sp12_h_r_17')
// (28, 31, 'sp12_h_r_18')
// (29, 31, 'sp12_h_r_21')
// (30, 31, 'sp12_h_r_22')
// (31, 31, 'sp12_h_l_22')
// (31, 31, 'sp12_v_t_22')
// (31, 32, 'sp12_v_b_22')
// (31, 33, 'io_1/OUT_ENB')
// (31, 33, 'local_g1_5')
// (31, 33, 'span12_vert_21')

reg n1380 = 0;
// (18, 19, 'neigh_op_tnr_4')
// (18, 20, 'neigh_op_rgt_4')
// (18, 21, 'neigh_op_bnr_4')
// (19, 19, 'neigh_op_top_4')
// (19, 20, 'local_g1_4')
// (19, 20, 'lutff_4/in_1')
// (19, 20, 'lutff_4/out')
// (19, 20, 'sp12_h_r_0')
// (19, 21, 'neigh_op_bot_4')
// (20, 19, 'neigh_op_tnl_4')
// (20, 20, 'neigh_op_lft_4')
// (20, 20, 'sp12_h_r_3')
// (20, 21, 'neigh_op_bnl_4')
// (21, 20, 'sp12_h_r_4')
// (22, 20, 'sp12_h_r_7')
// (23, 20, 'sp12_h_r_8')
// (24, 20, 'sp12_h_r_11')
// (25, 20, 'sp12_h_r_12')
// (26, 20, 'sp12_h_r_15')
// (27, 20, 'sp12_h_r_16')
// (27, 33, 'span4_horz_r_2')
// (28, 20, 'sp12_h_r_19')
// (28, 33, 'span4_horz_r_6')
// (29, 20, 'sp12_h_r_20')
// (29, 33, 'io_0/OUT_ENB')
// (29, 33, 'local_g1_2')
// (29, 33, 'span4_horz_r_10')
// (30, 20, 'sp12_h_r_23')
// (30, 29, 'sp4_r_v_b_37')
// (30, 30, 'sp4_r_v_b_24')
// (30, 31, 'sp4_r_v_b_13')
// (30, 32, 'sp4_r_v_b_0')
// (30, 33, 'span4_horz_r_14')
// (31, 20, 'sp12_h_l_23')
// (31, 20, 'sp12_v_t_23')
// (31, 21, 'sp12_v_b_23')
// (31, 22, 'sp12_v_b_20')
// (31, 23, 'sp12_v_b_19')
// (31, 24, 'sp12_v_b_16')
// (31, 25, 'sp12_v_b_15')
// (31, 26, 'sp12_v_b_12')
// (31, 27, 'sp12_v_b_11')
// (31, 28, 'sp12_v_b_8')
// (31, 28, 'sp4_v_t_37')
// (31, 29, 'sp12_v_b_7')
// (31, 29, 'sp4_v_b_37')
// (31, 30, 'sp12_v_b_4')
// (31, 30, 'sp4_v_b_24')
// (31, 31, 'sp12_v_b_3')
// (31, 31, 'sp4_v_b_13')
// (31, 32, 'sp12_v_b_0')
// (31, 32, 'sp4_v_b_0')
// (31, 32, 'sp4_v_t_37')
// (31, 33, 'span4_horz_l_14')
// (31, 33, 'span4_vert_37')

wire n1381;
// (18, 19, 'sp12_h_r_0')
// (18, 20, 'sp4_r_v_b_38')
// (18, 21, 'sp4_r_v_b_27')
// (18, 22, 'sp4_r_v_b_14')
// (18, 23, 'sp4_r_v_b_3')
// (19, 19, 'sp12_h_r_3')
// (19, 19, 'sp4_h_r_3')
// (19, 19, 'sp4_v_t_38')
// (19, 20, 'sp4_v_b_38')
// (19, 21, 'local_g2_3')
// (19, 21, 'lutff_5/in_2')
// (19, 21, 'sp4_v_b_27')
// (19, 22, 'sp4_v_b_14')
// (19, 23, 'sp4_v_b_3')
// (20, 19, 'sp12_h_r_4')
// (20, 19, 'sp4_h_r_14')
// (21, 19, 'sp12_h_r_7')
// (21, 19, 'sp4_h_r_27')
// (22, 19, 'sp12_h_r_8')
// (22, 19, 'sp4_h_r_38')
// (23, 19, 'sp12_h_r_11')
// (23, 19, 'sp4_h_l_38')
// (24, 19, 'sp12_h_r_12')
// (25, 19, 'sp12_h_r_15')
// (26, 19, 'sp12_h_r_16')
// (27, 19, 'sp12_h_r_19')
// (28, 19, 'sp12_h_r_20')
// (29, 19, 'sp12_h_r_23')
// (29, 32, 'neigh_op_tnr_2')
// (29, 32, 'neigh_op_tnr_6')
// (30, 19, 'sp12_h_l_23')
// (30, 19, 'sp12_v_t_23')
// (30, 20, 'sp12_v_b_23')
// (30, 21, 'sp12_v_b_20')
// (30, 22, 'sp12_v_b_19')
// (30, 23, 'sp12_v_b_16')
// (30, 24, 'sp12_v_b_15')
// (30, 25, 'sp12_v_b_12')
// (30, 26, 'sp12_v_b_11')
// (30, 27, 'sp12_v_b_8')
// (30, 28, 'sp12_v_b_7')
// (30, 29, 'sp12_v_b_4')
// (30, 30, 'sp12_v_b_3')
// (30, 31, 'sp12_v_b_0')
// (30, 31, 'sp12_v_t_23')
// (30, 32, 'neigh_op_top_2')
// (30, 32, 'neigh_op_top_6')
// (30, 32, 'sp12_v_b_23')
// (30, 33, 'io_1/D_IN_0')
// (30, 33, 'span12_vert_20')
// (31, 32, 'neigh_op_tnl_2')
// (31, 32, 'neigh_op_tnl_6')

wire n1382;
// (18, 19, 'sp4_r_v_b_44')
// (18, 20, 'sp4_r_v_b_33')
// (18, 21, 'sp4_r_v_b_20')
// (18, 22, 'sp4_r_v_b_9')
// (19, 18, 'sp4_h_r_9')
// (19, 18, 'sp4_v_t_44')
// (19, 19, 'sp4_v_b_44')
// (19, 20, 'sp4_v_b_33')
// (19, 21, 'local_g1_4')
// (19, 21, 'lutff_3/in_2')
// (19, 21, 'sp4_v_b_20')
// (19, 22, 'sp4_v_b_9')
// (20, 18, 'sp4_h_r_20')
// (21, 18, 'sp4_h_r_33')
// (22, 14, 'sp12_h_r_0')
// (22, 15, 'sp4_r_v_b_44')
// (22, 16, 'sp4_r_v_b_33')
// (22, 17, 'sp4_r_v_b_20')
// (22, 18, 'sp4_h_r_44')
// (22, 18, 'sp4_r_v_b_9')
// (23, 14, 'sp12_h_r_3')
// (23, 14, 'sp4_h_r_3')
// (23, 14, 'sp4_v_t_44')
// (23, 15, 'sp4_v_b_44')
// (23, 16, 'sp4_v_b_33')
// (23, 17, 'sp4_v_b_20')
// (23, 18, 'sp4_h_l_44')
// (23, 18, 'sp4_v_b_9')
// (24, 14, 'sp12_h_r_4')
// (24, 14, 'sp4_h_r_14')
// (25, 14, 'sp12_h_r_7')
// (25, 14, 'sp4_h_r_27')
// (26, 14, 'sp12_h_r_8')
// (26, 14, 'sp4_h_r_38')
// (27, 14, 'sp12_h_r_11')
// (27, 14, 'sp4_h_l_38')
// (28, 14, 'sp12_h_r_12')
// (29, 14, 'sp12_h_r_15')
// (30, 14, 'sp12_h_r_16')
// (31, 14, 'sp12_h_r_19')
// (32, 13, 'neigh_op_tnr_2')
// (32, 13, 'neigh_op_tnr_6')
// (32, 14, 'neigh_op_rgt_2')
// (32, 14, 'neigh_op_rgt_6')
// (32, 14, 'sp12_h_r_20')
// (32, 15, 'neigh_op_bnr_2')
// (32, 15, 'neigh_op_bnr_6')
// (33, 14, 'io_1/D_IN_0')
// (33, 14, 'span12_horz_20')

reg n1383 = 0;
// (18, 20, 'local_g0_3')
// (18, 20, 'lutff_4/in_1')
// (18, 20, 'sp4_h_r_11')
// (19, 20, 'sp4_h_r_22')
// (20, 20, 'sp4_h_r_35')
// (21, 20, 'neigh_op_tnr_4')
// (21, 20, 'sp4_h_r_46')
// (21, 21, 'neigh_op_rgt_4')
// (21, 21, 'sp4_r_v_b_40')
// (21, 22, 'neigh_op_bnr_4')
// (21, 22, 'sp4_r_v_b_29')
// (21, 23, 'sp4_r_v_b_16')
// (21, 24, 'sp4_r_v_b_5')
// (22, 20, 'neigh_op_top_4')
// (22, 20, 'sp4_h_l_46')
// (22, 20, 'sp4_v_t_40')
// (22, 21, 'lutff_4/out')
// (22, 21, 'sp4_v_b_40')
// (22, 22, 'neigh_op_bot_4')
// (22, 22, 'sp4_v_b_29')
// (22, 23, 'sp4_v_b_16')
// (22, 24, 'sp4_v_b_5')
// (23, 20, 'neigh_op_tnl_4')
// (23, 21, 'neigh_op_lft_4')
// (23, 22, 'neigh_op_bnl_4')

reg n1384 = 0;
// (18, 20, 'local_g1_0')
// (18, 20, 'lutff_0/in_1')
// (18, 20, 'sp4_h_r_0')
// (19, 19, 'neigh_op_tnr_4')
// (19, 20, 'neigh_op_rgt_4')
// (19, 20, 'sp4_h_r_13')
// (19, 21, 'neigh_op_bnr_4')
// (20, 19, 'neigh_op_top_4')
// (20, 20, 'lutff_4/out')
// (20, 20, 'sp4_h_r_24')
// (20, 21, 'neigh_op_bot_4')
// (21, 19, 'neigh_op_tnl_4')
// (21, 20, 'neigh_op_lft_4')
// (21, 20, 'sp4_h_r_37')
// (21, 21, 'neigh_op_bnl_4')
// (22, 20, 'sp4_h_l_37')

wire n1385;
// (18, 20, 'lutff_0/lout')
// (18, 20, 'lutff_1/in_2')

wire n1386;
// (18, 20, 'lutff_1/lout')
// (18, 20, 'lutff_2/in_2')

reg n1387 = 0;
// (18, 20, 'sp12_h_r_1')
// (18, 20, 'sp12_v_t_22')
// (18, 21, 'sp12_v_b_22')
// (18, 22, 'sp12_v_b_21')
// (18, 23, 'sp12_v_b_18')
// (18, 24, 'sp12_v_b_17')
// (18, 25, 'local_g3_6')
// (18, 25, 'lutff_4/in_1')
// (18, 25, 'sp12_v_b_14')
// (18, 26, 'sp12_v_b_13')
// (18, 27, 'sp12_v_b_10')
// (18, 28, 'sp12_v_b_9')
// (18, 29, 'sp12_v_b_6')
// (18, 30, 'sp12_v_b_5')
// (18, 31, 'sp12_v_b_2')
// (18, 32, 'sp12_v_b_1')
// (19, 20, 'sp12_h_r_2')
// (20, 19, 'neigh_op_tnr_7')
// (20, 20, 'neigh_op_rgt_7')
// (20, 20, 'sp12_h_r_5')
// (20, 21, 'neigh_op_bnr_7')
// (21, 19, 'neigh_op_top_7')
// (21, 20, 'lutff_7/out')
// (21, 20, 'sp12_h_r_6')
// (21, 21, 'neigh_op_bot_7')
// (22, 19, 'neigh_op_tnl_7')
// (22, 20, 'neigh_op_lft_7')
// (22, 20, 'sp12_h_r_9')
// (22, 21, 'neigh_op_bnl_7')
// (23, 20, 'sp12_h_r_10')
// (24, 20, 'sp12_h_r_13')
// (25, 20, 'sp12_h_r_14')
// (26, 20, 'sp12_h_r_17')
// (27, 20, 'sp12_h_r_18')
// (28, 20, 'sp12_h_r_21')
// (29, 20, 'sp12_h_r_22')
// (30, 20, 'sp12_h_l_22')

wire n1388;
// (18, 20, 'sp4_r_v_b_37')
// (18, 21, 'sp4_r_v_b_24')
// (18, 22, 'sp4_r_v_b_13')
// (18, 23, 'sp4_r_v_b_0')
// (19, 19, 'sp4_h_r_0')
// (19, 19, 'sp4_v_t_37')
// (19, 20, 'sp4_v_b_37')
// (19, 21, 'local_g2_0')
// (19, 21, 'lutff_4/in_0')
// (19, 21, 'sp4_v_b_24')
// (19, 22, 'sp4_v_b_13')
// (19, 23, 'sp4_v_b_0')
// (20, 19, 'sp4_h_r_13')
// (21, 19, 'sp4_h_r_24')
// (22, 16, 'sp4_r_v_b_42')
// (22, 17, 'sp4_r_v_b_31')
// (22, 18, 'sp4_r_v_b_18')
// (22, 19, 'sp4_h_r_37')
// (22, 19, 'sp4_r_v_b_7')
// (23, 15, 'sp4_h_r_1')
// (23, 15, 'sp4_v_t_42')
// (23, 16, 'sp4_v_b_42')
// (23, 17, 'sp4_v_b_31')
// (23, 18, 'sp4_v_b_18')
// (23, 19, 'sp4_h_l_37')
// (23, 19, 'sp4_v_b_7')
// (24, 15, 'sp12_h_r_0')
// (24, 15, 'sp4_h_r_12')
// (25, 15, 'sp12_h_r_3')
// (25, 15, 'sp4_h_r_25')
// (26, 15, 'sp12_h_r_4')
// (26, 15, 'sp4_h_r_36')
// (27, 15, 'sp12_h_r_7')
// (27, 15, 'sp4_h_l_36')
// (28, 15, 'sp12_h_r_8')
// (29, 15, 'sp12_h_r_11')
// (30, 15, 'sp12_h_r_12')
// (31, 15, 'sp12_h_r_15')
// (32, 14, 'neigh_op_tnr_0')
// (32, 14, 'neigh_op_tnr_4')
// (32, 15, 'neigh_op_rgt_0')
// (32, 15, 'neigh_op_rgt_4')
// (32, 15, 'sp12_h_r_16')
// (32, 16, 'neigh_op_bnr_0')
// (32, 16, 'neigh_op_bnr_4')
// (33, 15, 'io_0/D_IN_0')
// (33, 15, 'span12_horz_16')

reg n1389 = 0;
// (18, 21, 'neigh_op_tnr_0')
// (18, 22, 'neigh_op_rgt_0')
// (18, 23, 'neigh_op_bnr_0')
// (19, 21, 'neigh_op_top_0')
// (19, 22, 'local_g3_0')
// (19, 22, 'lutff_0/in_1')
// (19, 22, 'lutff_0/out')
// (19, 23, 'neigh_op_bot_0')
// (20, 21, 'neigh_op_tnl_0')
// (20, 22, 'local_g0_0')
// (20, 22, 'lutff_0/in_0')
// (20, 22, 'neigh_op_lft_0')
// (20, 23, 'neigh_op_bnl_0')

reg n1390 = 0;
// (18, 21, 'neigh_op_tnr_1')
// (18, 22, 'neigh_op_rgt_1')
// (18, 23, 'neigh_op_bnr_1')
// (19, 21, 'neigh_op_top_1')
// (19, 22, 'local_g3_1')
// (19, 22, 'lutff_1/in_1')
// (19, 22, 'lutff_1/out')
// (19, 23, 'neigh_op_bot_1')
// (20, 21, 'neigh_op_tnl_1')
// (20, 22, 'local_g0_1')
// (20, 22, 'lutff_4/in_1')
// (20, 22, 'neigh_op_lft_1')
// (20, 23, 'neigh_op_bnl_1')

reg n1391 = 0;
// (18, 21, 'neigh_op_tnr_2')
// (18, 22, 'neigh_op_rgt_2')
// (18, 23, 'neigh_op_bnr_2')
// (19, 21, 'neigh_op_top_2')
// (19, 22, 'local_g1_2')
// (19, 22, 'lutff_2/in_1')
// (19, 22, 'lutff_2/out')
// (19, 22, 'sp4_h_r_4')
// (19, 23, 'neigh_op_bot_2')
// (20, 21, 'neigh_op_tnl_2')
// (20, 22, 'local_g1_1')
// (20, 22, 'lutff_4/in_0')
// (20, 22, 'neigh_op_lft_2')
// (20, 22, 'sp4_h_r_17')
// (20, 23, 'neigh_op_bnl_2')
// (21, 22, 'sp4_h_r_28')
// (22, 22, 'sp4_h_r_41')
// (23, 22, 'sp4_h_l_41')

reg n1392 = 0;
// (18, 21, 'neigh_op_tnr_3')
// (18, 22, 'neigh_op_rgt_3')
// (18, 23, 'neigh_op_bnr_3')
// (19, 21, 'neigh_op_top_3')
// (19, 22, 'local_g3_3')
// (19, 22, 'lutff_3/in_1')
// (19, 22, 'lutff_3/out')
// (19, 23, 'neigh_op_bot_3')
// (20, 21, 'neigh_op_tnl_3')
// (20, 22, 'local_g1_3')
// (20, 22, 'lutff_3/in_3')
// (20, 22, 'neigh_op_lft_3')
// (20, 23, 'neigh_op_bnl_3')

reg n1393 = 0;
// (18, 21, 'neigh_op_tnr_4')
// (18, 22, 'neigh_op_rgt_4')
// (18, 23, 'neigh_op_bnr_4')
// (19, 21, 'neigh_op_top_4')
// (19, 22, 'local_g3_4')
// (19, 22, 'lutff_4/in_1')
// (19, 22, 'lutff_4/out')
// (19, 23, 'neigh_op_bot_4')
// (20, 21, 'neigh_op_tnl_4')
// (20, 22, 'local_g0_4')
// (20, 22, 'lutff_0/in_2')
// (20, 22, 'neigh_op_lft_4')
// (20, 23, 'neigh_op_bnl_4')

reg n1394 = 0;
// (18, 21, 'neigh_op_tnr_5')
// (18, 22, 'neigh_op_rgt_5')
// (18, 23, 'neigh_op_bnr_5')
// (19, 21, 'neigh_op_top_5')
// (19, 22, 'local_g1_5')
// (19, 22, 'lutff_5/in_1')
// (19, 22, 'lutff_5/out')
// (19, 23, 'neigh_op_bot_5')
// (20, 21, 'neigh_op_tnl_5')
// (20, 22, 'local_g0_5')
// (20, 22, 'lutff_0/in_3')
// (20, 22, 'neigh_op_lft_5')
// (20, 23, 'neigh_op_bnl_5')

reg n1395 = 0;
// (18, 21, 'neigh_op_tnr_6')
// (18, 22, 'neigh_op_rgt_6')
// (18, 23, 'neigh_op_bnr_6')
// (19, 21, 'neigh_op_top_6')
// (19, 22, 'local_g1_6')
// (19, 22, 'lutff_6/in_1')
// (19, 22, 'lutff_6/out')
// (19, 23, 'neigh_op_bot_6')
// (20, 21, 'neigh_op_tnl_6')
// (20, 22, 'local_g0_6')
// (20, 22, 'lutff_3/in_1')
// (20, 22, 'neigh_op_lft_6')
// (20, 23, 'neigh_op_bnl_6')

reg n1396 = 0;
// (18, 21, 'neigh_op_tnr_7')
// (18, 22, 'neigh_op_rgt_7')
// (18, 23, 'neigh_op_bnr_7')
// (19, 21, 'neigh_op_top_7')
// (19, 22, 'local_g1_7')
// (19, 22, 'lutff_7/in_1')
// (19, 22, 'lutff_7/out')
// (19, 23, 'neigh_op_bot_7')
// (20, 21, 'neigh_op_tnl_7')
// (20, 22, 'local_g0_7')
// (20, 22, 'lutff_0/in_1')
// (20, 22, 'neigh_op_lft_7')
// (20, 23, 'neigh_op_bnl_7')

wire n1397;
// (18, 21, 'sp4_r_v_b_39')
// (18, 22, 'sp4_r_v_b_26')
// (18, 23, 'sp4_r_v_b_15')
// (18, 24, 'sp4_r_v_b_2')
// (19, 20, 'sp4_h_r_8')
// (19, 20, 'sp4_v_t_39')
// (19, 21, 'local_g3_7')
// (19, 21, 'lutff_7/in_1')
// (19, 21, 'sp4_v_b_39')
// (19, 22, 'sp4_v_b_26')
// (19, 23, 'sp4_v_b_15')
// (19, 24, 'sp4_v_b_2')
// (20, 20, 'sp4_h_r_21')
// (21, 20, 'sp4_h_r_32')
// (22, 16, 'sp12_h_r_0')
// (22, 17, 'sp4_r_v_b_38')
// (22, 18, 'sp4_r_v_b_27')
// (22, 19, 'sp4_r_v_b_14')
// (22, 20, 'sp4_h_r_45')
// (22, 20, 'sp4_r_v_b_3')
// (23, 16, 'sp12_h_r_3')
// (23, 16, 'sp4_h_r_3')
// (23, 16, 'sp4_v_t_38')
// (23, 17, 'sp4_v_b_38')
// (23, 18, 'sp4_v_b_27')
// (23, 19, 'sp4_v_b_14')
// (23, 20, 'sp4_h_l_45')
// (23, 20, 'sp4_v_b_3')
// (24, 16, 'sp12_h_r_4')
// (24, 16, 'sp4_h_r_14')
// (25, 16, 'sp12_h_r_7')
// (25, 16, 'sp4_h_r_27')
// (26, 16, 'sp12_h_r_8')
// (26, 16, 'sp4_h_r_38')
// (27, 16, 'sp12_h_r_11')
// (27, 16, 'sp4_h_l_38')
// (28, 16, 'sp12_h_r_12')
// (29, 16, 'sp12_h_r_15')
// (30, 16, 'sp12_h_r_16')
// (31, 16, 'sp12_h_r_19')
// (32, 15, 'neigh_op_tnr_2')
// (32, 15, 'neigh_op_tnr_6')
// (32, 16, 'neigh_op_rgt_2')
// (32, 16, 'neigh_op_rgt_6')
// (32, 16, 'sp12_h_r_20')
// (32, 17, 'neigh_op_bnr_2')
// (32, 17, 'neigh_op_bnr_6')
// (33, 16, 'io_1/D_IN_0')
// (33, 16, 'span12_horz_20')

wire n1398;
// (18, 21, 'sp4_r_v_b_42')
// (18, 22, 'sp4_r_v_b_31')
// (18, 23, 'sp4_r_v_b_18')
// (18, 24, 'sp4_r_v_b_7')
// (19, 20, 'sp4_h_r_1')
// (19, 20, 'sp4_v_t_42')
// (19, 21, 'local_g2_2')
// (19, 21, 'lutff_6/in_0')
// (19, 21, 'sp4_v_b_42')
// (19, 22, 'sp4_v_b_31')
// (19, 23, 'sp4_v_b_18')
// (19, 24, 'sp4_v_b_7')
// (20, 20, 'sp4_h_r_12')
// (21, 20, 'sp4_h_r_25')
// (22, 17, 'sp4_r_v_b_36')
// (22, 18, 'sp4_r_v_b_25')
// (22, 19, 'sp4_r_v_b_12')
// (22, 20, 'sp4_h_r_36')
// (22, 20, 'sp4_r_v_b_1')
// (23, 16, 'sp4_h_r_1')
// (23, 16, 'sp4_v_t_36')
// (23, 17, 'sp4_v_b_36')
// (23, 18, 'sp4_v_b_25')
// (23, 19, 'sp4_v_b_12')
// (23, 20, 'sp4_h_l_36')
// (23, 20, 'sp4_v_b_1')
// (24, 16, 'sp12_h_r_0')
// (24, 16, 'sp4_h_r_12')
// (25, 16, 'sp12_h_r_3')
// (25, 16, 'sp4_h_r_25')
// (26, 16, 'sp12_h_r_4')
// (26, 16, 'sp4_h_r_36')
// (27, 16, 'sp12_h_r_7')
// (27, 16, 'sp4_h_l_36')
// (28, 16, 'sp12_h_r_8')
// (29, 16, 'sp12_h_r_11')
// (30, 16, 'sp12_h_r_12')
// (31, 16, 'sp12_h_r_15')
// (32, 15, 'neigh_op_tnr_0')
// (32, 15, 'neigh_op_tnr_4')
// (32, 16, 'neigh_op_rgt_0')
// (32, 16, 'neigh_op_rgt_4')
// (32, 16, 'sp12_h_r_16')
// (32, 17, 'neigh_op_bnr_0')
// (32, 17, 'neigh_op_bnr_4')
// (33, 16, 'io_0/D_IN_0')
// (33, 16, 'span12_horz_16')

wire n1399;
// (18, 22, 'lutff_2/lout')
// (18, 22, 'lutff_3/in_2')

reg n1400 = 0;
// (18, 22, 'neigh_op_tnr_1')
// (18, 23, 'neigh_op_rgt_1')
// (18, 24, 'neigh_op_bnr_1')
// (19, 20, 'sp12_v_t_22')
// (19, 21, 'sp12_v_b_22')
// (19, 22, 'neigh_op_top_1')
// (19, 22, 'sp12_v_b_21')
// (19, 23, 'local_g0_1')
// (19, 23, 'lutff_1/in_2')
// (19, 23, 'lutff_1/out')
// (19, 23, 'sp12_v_b_18')
// (19, 24, 'neigh_op_bot_1')
// (19, 24, 'sp12_v_b_17')
// (19, 25, 'sp12_v_b_14')
// (19, 26, 'sp12_v_b_13')
// (19, 27, 'sp12_v_b_10')
// (19, 28, 'sp12_v_b_9')
// (19, 29, 'sp12_v_b_6')
// (19, 30, 'sp12_v_b_5')
// (19, 31, 'sp12_v_b_2')
// (19, 32, 'sp12_h_r_1')
// (19, 32, 'sp12_v_b_1')
// (20, 22, 'neigh_op_tnl_1')
// (20, 23, 'neigh_op_lft_1')
// (20, 24, 'neigh_op_bnl_1')
// (20, 32, 'sp12_h_r_2')
// (21, 32, 'sp12_h_r_5')
// (22, 32, 'sp12_h_r_6')
// (23, 32, 'sp12_h_r_9')
// (24, 32, 'sp12_h_r_10')
// (25, 32, 'sp12_h_r_13')
// (26, 32, 'sp12_h_r_14')
// (27, 32, 'sp12_h_r_17')
// (28, 32, 'sp12_h_r_18')
// (29, 32, 'sp12_h_r_21')
// (30, 32, 'sp12_h_r_22')
// (31, 32, 'sp12_h_l_22')
// (31, 32, 'sp12_v_t_22')
// (31, 33, 'io_0/OUT_ENB')
// (31, 33, 'local_g1_6')
// (31, 33, 'span12_vert_22')

reg n1401 = 0;
// (18, 22, 'neigh_op_tnr_3')
// (18, 23, 'neigh_op_rgt_3')
// (18, 24, 'neigh_op_bnr_3')
// (19, 10, 'sp12_h_r_1')
// (19, 10, 'sp12_v_t_22')
// (19, 11, 'sp12_v_b_22')
// (19, 12, 'sp12_v_b_21')
// (19, 13, 'sp12_v_b_18')
// (19, 14, 'sp12_v_b_17')
// (19, 15, 'sp12_v_b_14')
// (19, 16, 'sp12_v_b_13')
// (19, 17, 'sp12_v_b_10')
// (19, 18, 'sp12_v_b_9')
// (19, 19, 'sp12_v_b_6')
// (19, 20, 'sp12_v_b_5')
// (19, 21, 'sp12_v_b_2')
// (19, 22, 'neigh_op_top_3')
// (19, 22, 'sp12_v_b_1')
// (19, 22, 'sp12_v_t_22')
// (19, 23, 'local_g0_3')
// (19, 23, 'lutff_3/in_2')
// (19, 23, 'lutff_3/out')
// (19, 23, 'sp12_v_b_22')
// (19, 24, 'neigh_op_bot_3')
// (19, 24, 'sp12_v_b_21')
// (19, 25, 'sp12_v_b_18')
// (19, 26, 'sp12_v_b_17')
// (19, 27, 'sp12_v_b_14')
// (19, 28, 'sp12_v_b_13')
// (19, 29, 'sp12_v_b_10')
// (19, 30, 'sp12_v_b_9')
// (19, 31, 'sp12_v_b_6')
// (19, 32, 'sp12_v_b_5')
// (19, 33, 'span12_vert_2')
// (20, 10, 'sp12_h_r_2')
// (20, 22, 'neigh_op_tnl_3')
// (20, 23, 'neigh_op_lft_3')
// (20, 24, 'neigh_op_bnl_3')
// (21, 10, 'sp12_h_r_5')
// (22, 10, 'sp12_h_r_6')
// (23, 10, 'sp12_h_r_9')
// (24, 10, 'sp12_h_r_10')
// (25, 10, 'sp12_h_r_13')
// (26, 10, 'sp12_h_r_14')
// (27, 10, 'sp12_h_r_17')
// (28, 10, 'sp12_h_r_18')
// (29, 10, 'sp12_h_r_21')
// (29, 10, 'sp4_h_r_10')
// (30, 10, 'sp12_h_r_22')
// (30, 10, 'sp4_h_r_23')
// (31, 10, 'sp12_h_l_22')
// (31, 10, 'sp4_h_r_34')
// (32, 10, 'sp4_h_r_47')
// (33, 10, 'io_1/OUT_ENB')
// (33, 10, 'local_g1_7')
// (33, 10, 'span4_horz_47')

reg n1402 = 0;
// (18, 22, 'neigh_op_tnr_4')
// (18, 23, 'neigh_op_rgt_4')
// (18, 24, 'neigh_op_bnr_4')
// (19, 22, 'neigh_op_top_4')
// (19, 23, 'local_g0_4')
// (19, 23, 'lutff_4/in_0')
// (19, 23, 'lutff_4/out')
// (19, 23, 'sp12_h_r_0')
// (19, 24, 'neigh_op_bot_4')
// (20, 22, 'neigh_op_tnl_4')
// (20, 23, 'neigh_op_lft_4')
// (20, 23, 'sp12_h_r_3')
// (20, 24, 'neigh_op_bnl_4')
// (21, 23, 'sp12_h_r_4')
// (22, 23, 'sp12_h_r_7')
// (23, 23, 'sp12_h_r_8')
// (24, 23, 'sp12_h_r_11')
// (25, 23, 'sp12_h_r_12')
// (26, 23, 'sp12_h_r_15')
// (27, 23, 'sp12_h_r_16')
// (28, 23, 'sp12_h_r_19')
// (29, 23, 'sp12_h_r_20')
// (30, 23, 'sp12_h_r_23')
// (30, 23, 'sp4_h_r_1')
// (31, 23, 'sp12_h_l_23')
// (31, 23, 'sp12_h_r_0')
// (31, 23, 'sp4_h_r_12')
// (32, 23, 'sp12_h_r_3')
// (32, 23, 'sp4_h_r_25')
// (33, 15, 'span4_vert_t_12')
// (33, 16, 'io_0/OUT_ENB')
// (33, 16, 'local_g1_4')
// (33, 16, 'span4_vert_b_12')
// (33, 17, 'span4_vert_b_8')
// (33, 18, 'span4_vert_b_4')
// (33, 19, 'span4_vert_b_0')
// (33, 19, 'span4_vert_t_12')
// (33, 20, 'span4_vert_b_12')
// (33, 21, 'span4_vert_b_8')
// (33, 22, 'span4_vert_b_4')
// (33, 23, 'span12_horz_3')
// (33, 23, 'span4_horz_25')
// (33, 23, 'span4_vert_b_0')

reg n1403 = 0;
// (18, 22, 'neigh_op_tnr_5')
// (18, 23, 'neigh_op_rgt_5')
// (18, 23, 'sp12_h_r_1')
// (18, 24, 'neigh_op_bnr_5')
// (19, 22, 'neigh_op_top_5')
// (19, 23, 'local_g2_5')
// (19, 23, 'lutff_5/in_2')
// (19, 23, 'lutff_5/out')
// (19, 23, 'sp12_h_r_2')
// (19, 24, 'neigh_op_bot_5')
// (20, 22, 'neigh_op_tnl_5')
// (20, 23, 'neigh_op_lft_5')
// (20, 23, 'sp12_h_r_5')
// (20, 24, 'neigh_op_bnl_5')
// (21, 23, 'sp12_h_r_6')
// (22, 23, 'sp12_h_r_9')
// (22, 23, 'sp4_h_r_4')
// (23, 23, 'sp12_h_r_10')
// (23, 23, 'sp4_h_r_17')
// (24, 23, 'sp12_h_r_13')
// (24, 23, 'sp4_h_r_28')
// (25, 23, 'sp12_h_r_14')
// (25, 23, 'sp4_h_r_41')
// (25, 24, 'sp4_r_v_b_44')
// (25, 25, 'sp4_r_v_b_33')
// (25, 26, 'sp4_r_v_b_20')
// (25, 27, 'sp4_r_v_b_9')
// (25, 28, 'sp4_r_v_b_40')
// (25, 29, 'sp4_r_v_b_29')
// (25, 30, 'sp4_r_v_b_16')
// (25, 31, 'sp4_r_v_b_5')
// (25, 32, 'sp4_r_v_b_36')
// (26, 23, 'sp12_h_r_17')
// (26, 23, 'sp4_h_l_41')
// (26, 23, 'sp4_v_t_44')
// (26, 24, 'sp4_v_b_44')
// (26, 25, 'sp4_v_b_33')
// (26, 26, 'sp4_v_b_20')
// (26, 27, 'sp4_v_b_9')
// (26, 27, 'sp4_v_t_40')
// (26, 28, 'sp4_v_b_40')
// (26, 29, 'sp4_v_b_29')
// (26, 30, 'sp4_v_b_16')
// (26, 31, 'sp4_v_b_5')
// (26, 31, 'sp4_v_t_36')
// (26, 32, 'sp4_v_b_36')
// (26, 33, 'span4_horz_r_0')
// (26, 33, 'span4_vert_25')
// (27, 23, 'sp12_h_r_18')
// (27, 33, 'span4_horz_r_4')
// (28, 23, 'sp12_h_r_21')
// (28, 33, 'span4_horz_r_8')
// (29, 23, 'sp12_h_r_22')
// (29, 33, 'io_1/OUT_ENB')
// (29, 33, 'local_g0_4')
// (29, 33, 'span4_horz_r_12')
// (30, 23, 'sp12_h_l_22')
// (30, 33, 'span4_horz_l_12')

reg n1404 = 0;
// (18, 22, 'neigh_op_tnr_6')
// (18, 23, 'neigh_op_rgt_6')
// (18, 24, 'neigh_op_bnr_6')
// (19, 17, 'sp12_v_t_23')
// (19, 18, 'sp12_v_b_23')
// (19, 19, 'sp12_v_b_20')
// (19, 20, 'sp12_v_b_19')
// (19, 21, 'sp12_v_b_16')
// (19, 22, 'neigh_op_top_6')
// (19, 22, 'sp12_v_b_15')
// (19, 23, 'local_g2_6')
// (19, 23, 'lutff_6/in_0')
// (19, 23, 'lutff_6/out')
// (19, 23, 'sp12_v_b_12')
// (19, 24, 'neigh_op_bot_6')
// (19, 24, 'sp12_v_b_11')
// (19, 25, 'sp12_v_b_8')
// (19, 26, 'sp12_v_b_7')
// (19, 27, 'sp12_v_b_4')
// (19, 28, 'sp12_v_b_3')
// (19, 29, 'sp12_h_r_0')
// (19, 29, 'sp12_v_b_0')
// (20, 22, 'neigh_op_tnl_6')
// (20, 23, 'neigh_op_lft_6')
// (20, 24, 'neigh_op_bnl_6')
// (20, 29, 'sp12_h_r_3')
// (21, 29, 'sp12_h_r_4')
// (22, 29, 'sp12_h_r_7')
// (23, 29, 'sp12_h_r_8')
// (24, 29, 'sp12_h_r_11')
// (24, 29, 'sp4_h_r_7')
// (25, 29, 'sp12_h_r_12')
// (25, 29, 'sp4_h_r_18')
// (26, 29, 'sp12_h_r_15')
// (26, 29, 'sp4_h_r_31')
// (27, 29, 'sp12_h_r_16')
// (27, 29, 'sp4_h_r_42')
// (27, 30, 'sp4_r_v_b_37')
// (27, 31, 'sp4_r_v_b_24')
// (27, 32, 'sp4_r_v_b_13')
// (28, 29, 'sp12_h_r_19')
// (28, 29, 'sp4_h_l_42')
// (28, 29, 'sp4_v_t_37')
// (28, 30, 'sp4_v_b_37')
// (28, 31, 'sp4_v_b_24')
// (28, 32, 'sp4_v_b_13')
// (28, 33, 'io_1/OUT_ENB')
// (28, 33, 'local_g0_0')
// (28, 33, 'span4_vert_0')
// (29, 29, 'sp12_h_r_20')
// (30, 29, 'sp12_h_r_23')
// (31, 29, 'sp12_h_l_23')

reg n1405 = 0;
// (18, 23, 'neigh_op_tnr_0')
// (18, 24, 'neigh_op_rgt_0')
// (18, 25, 'neigh_op_bnr_0')
// (19, 23, 'neigh_op_top_0')
// (19, 24, 'local_g3_0')
// (19, 24, 'lutff_0/in_1')
// (19, 24, 'lutff_0/out')
// (19, 25, 'neigh_op_bot_0')
// (20, 23, 'neigh_op_tnl_0')
// (20, 24, 'local_g0_0')
// (20, 24, 'lutff_1/in_1')
// (20, 24, 'neigh_op_lft_0')
// (20, 25, 'neigh_op_bnl_0')

reg n1406 = 0;
// (18, 23, 'neigh_op_tnr_1')
// (18, 24, 'neigh_op_rgt_1')
// (18, 25, 'neigh_op_bnr_1')
// (19, 23, 'neigh_op_top_1')
// (19, 24, 'local_g3_1')
// (19, 24, 'lutff_1/in_1')
// (19, 24, 'lutff_1/out')
// (19, 25, 'neigh_op_bot_1')
// (20, 23, 'neigh_op_tnl_1')
// (20, 24, 'local_g0_1')
// (20, 24, 'lutff_1/in_2')
// (20, 24, 'neigh_op_lft_1')
// (20, 25, 'neigh_op_bnl_1')

reg n1407 = 0;
// (18, 23, 'neigh_op_tnr_2')
// (18, 24, 'neigh_op_rgt_2')
// (18, 25, 'neigh_op_bnr_2')
// (19, 23, 'neigh_op_top_2')
// (19, 24, 'local_g1_2')
// (19, 24, 'lutff_2/in_1')
// (19, 24, 'lutff_2/out')
// (19, 25, 'neigh_op_bot_2')
// (20, 23, 'neigh_op_tnl_2')
// (20, 24, 'local_g1_2')
// (20, 24, 'lutff_2/in_3')
// (20, 24, 'neigh_op_lft_2')
// (20, 25, 'neigh_op_bnl_2')

reg n1408 = 0;
// (18, 23, 'neigh_op_tnr_3')
// (18, 24, 'neigh_op_rgt_3')
// (18, 25, 'neigh_op_bnr_3')
// (19, 23, 'neigh_op_top_3')
// (19, 24, 'local_g1_3')
// (19, 24, 'lutff_3/in_1')
// (19, 24, 'lutff_3/out')
// (19, 25, 'neigh_op_bot_3')
// (20, 23, 'neigh_op_tnl_3')
// (20, 24, 'local_g0_3')
// (20, 24, 'lutff_2/in_1')
// (20, 24, 'neigh_op_lft_3')
// (20, 25, 'neigh_op_bnl_3')

reg n1409 = 0;
// (18, 23, 'neigh_op_tnr_4')
// (18, 24, 'neigh_op_rgt_4')
// (18, 25, 'neigh_op_bnr_4')
// (19, 23, 'neigh_op_top_4')
// (19, 24, 'local_g3_4')
// (19, 24, 'lutff_4/in_1')
// (19, 24, 'lutff_4/out')
// (19, 25, 'neigh_op_bot_4')
// (20, 23, 'neigh_op_tnl_4')
// (20, 24, 'local_g0_4')
// (20, 24, 'lutff_7/in_3')
// (20, 24, 'neigh_op_lft_4')
// (20, 25, 'neigh_op_bnl_4')

reg n1410 = 0;
// (18, 23, 'neigh_op_tnr_5')
// (18, 24, 'neigh_op_rgt_5')
// (18, 25, 'neigh_op_bnr_5')
// (19, 23, 'neigh_op_top_5')
// (19, 24, 'local_g1_5')
// (19, 24, 'lutff_5/in_1')
// (19, 24, 'lutff_5/out')
// (19, 25, 'neigh_op_bot_5')
// (20, 23, 'neigh_op_tnl_5')
// (20, 24, 'local_g0_5')
// (20, 24, 'lutff_7/in_0')
// (20, 24, 'neigh_op_lft_5')
// (20, 25, 'neigh_op_bnl_5')

reg n1411 = 0;
// (18, 23, 'sp4_r_v_b_44')
// (18, 24, 'neigh_op_tnr_2')
// (18, 24, 'sp4_r_v_b_33')
// (18, 25, 'neigh_op_rgt_2')
// (18, 25, 'sp4_r_v_b_20')
// (18, 26, 'neigh_op_bnr_2')
// (18, 26, 'sp4_r_v_b_9')
// (19, 22, 'sp4_h_r_9')
// (19, 22, 'sp4_v_t_44')
// (19, 23, 'sp4_v_b_44')
// (19, 24, 'neigh_op_top_2')
// (19, 24, 'sp4_v_b_33')
// (19, 25, 'lutff_2/out')
// (19, 25, 'sp4_v_b_20')
// (19, 26, 'neigh_op_bot_2')
// (19, 26, 'sp4_v_b_9')
// (20, 22, 'sp4_h_r_20')
// (20, 24, 'neigh_op_tnl_2')
// (20, 25, 'neigh_op_lft_2')
// (20, 26, 'neigh_op_bnl_2')
// (21, 22, 'local_g3_1')
// (21, 22, 'lutff_3/in_3')
// (21, 22, 'sp4_h_r_33')
// (22, 22, 'sp4_h_r_44')
// (23, 22, 'sp4_h_l_44')

reg n1412 = 0;
// (18, 24, 'local_g1_4')
// (18, 24, 'lutff_2/in_1')
// (18, 24, 'sp4_h_r_4')
// (19, 24, 'sp4_h_r_17')
// (20, 24, 'sp4_h_r_28')
// (21, 17, 'sp4_r_v_b_38')
// (21, 18, 'sp4_r_v_b_27')
// (21, 19, 'sp4_r_v_b_14')
// (21, 20, 'sp4_r_v_b_3')
// (21, 21, 'sp4_r_v_b_46')
// (21, 22, 'sp4_r_v_b_35')
// (21, 23, 'sp4_r_v_b_22')
// (21, 24, 'sp4_h_r_41')
// (21, 24, 'sp4_r_v_b_11')
// (22, 15, 'neigh_op_tnr_7')
// (22, 16, 'neigh_op_rgt_7')
// (22, 16, 'sp4_h_r_3')
// (22, 16, 'sp4_v_t_38')
// (22, 17, 'neigh_op_bnr_7')
// (22, 17, 'sp4_v_b_38')
// (22, 18, 'sp4_v_b_27')
// (22, 19, 'sp4_v_b_14')
// (22, 20, 'sp4_v_b_3')
// (22, 20, 'sp4_v_t_46')
// (22, 21, 'sp4_v_b_46')
// (22, 22, 'sp4_v_b_35')
// (22, 23, 'sp4_v_b_22')
// (22, 24, 'sp4_h_l_41')
// (22, 24, 'sp4_v_b_11')
// (23, 15, 'neigh_op_top_7')
// (23, 16, 'lutff_7/out')
// (23, 16, 'sp4_h_r_14')
// (23, 17, 'neigh_op_bot_7')
// (24, 15, 'neigh_op_tnl_7')
// (24, 16, 'neigh_op_lft_7')
// (24, 16, 'sp4_h_r_27')
// (24, 17, 'neigh_op_bnl_7')
// (25, 16, 'sp4_h_r_38')
// (26, 16, 'sp4_h_l_38')

wire n1413;
// (18, 24, 'lutff_3/lout')
// (18, 24, 'lutff_4/in_2')

wire n1414;
// (18, 24, 'lutff_4/lout')
// (18, 24, 'lutff_5/in_2')

reg n1415 = 0;
// (18, 25, 'local_g0_2')
// (18, 25, 'lutff_6/in_0')
// (18, 25, 'sp4_h_r_10')
// (19, 24, 'neigh_op_tnr_1')
// (19, 25, 'neigh_op_rgt_1')
// (19, 25, 'sp4_h_r_23')
// (19, 26, 'neigh_op_bnr_1')
// (20, 24, 'neigh_op_top_1')
// (20, 25, 'lutff_1/out')
// (20, 25, 'sp4_h_r_34')
// (20, 26, 'neigh_op_bot_1')
// (21, 24, 'neigh_op_tnl_1')
// (21, 25, 'neigh_op_lft_1')
// (21, 25, 'sp4_h_r_47')
// (21, 26, 'neigh_op_bnl_1')
// (22, 25, 'sp4_h_l_47')

reg n1416 = 0;
// (18, 25, 'local_g0_3')
// (18, 25, 'lutff_6/in_3')
// (18, 25, 'sp4_h_r_3')
// (19, 25, 'sp4_h_r_14')
// (20, 25, 'sp4_h_r_27')
// (21, 22, 'neigh_op_tnr_1')
// (21, 22, 'sp4_r_v_b_47')
// (21, 23, 'neigh_op_rgt_1')
// (21, 23, 'sp4_r_v_b_34')
// (21, 24, 'neigh_op_bnr_1')
// (21, 24, 'sp4_r_v_b_23')
// (21, 25, 'sp4_h_r_38')
// (21, 25, 'sp4_r_v_b_10')
// (22, 21, 'sp4_v_t_47')
// (22, 22, 'neigh_op_top_1')
// (22, 22, 'sp4_v_b_47')
// (22, 23, 'lutff_1/out')
// (22, 23, 'sp4_v_b_34')
// (22, 24, 'neigh_op_bot_1')
// (22, 24, 'sp4_v_b_23')
// (22, 25, 'sp4_h_l_38')
// (22, 25, 'sp4_v_b_10')
// (23, 22, 'neigh_op_tnl_1')
// (23, 23, 'neigh_op_lft_1')
// (23, 24, 'neigh_op_bnl_1')

reg n1417 = 0;
// (18, 25, 'local_g0_7')
// (18, 25, 'lutff_4/in_3')
// (18, 25, 'sp4_h_r_7')
// (19, 25, 'sp4_h_r_18')
// (20, 25, 'sp4_h_r_31')
// (21, 22, 'sp4_r_v_b_42')
// (21, 23, 'neigh_op_tnr_1')
// (21, 23, 'sp4_r_v_b_31')
// (21, 24, 'neigh_op_rgt_1')
// (21, 24, 'sp4_r_v_b_18')
// (21, 25, 'neigh_op_bnr_1')
// (21, 25, 'sp4_h_r_42')
// (21, 25, 'sp4_r_v_b_7')
// (22, 21, 'sp4_v_t_42')
// (22, 22, 'sp4_v_b_42')
// (22, 23, 'neigh_op_top_1')
// (22, 23, 'sp4_v_b_31')
// (22, 24, 'lutff_1/out')
// (22, 24, 'sp4_v_b_18')
// (22, 25, 'neigh_op_bot_1')
// (22, 25, 'sp4_h_l_42')
// (22, 25, 'sp4_v_b_7')
// (23, 23, 'neigh_op_tnl_1')
// (23, 24, 'neigh_op_lft_1')
// (23, 25, 'neigh_op_bnl_1')

reg n1418 = 0;
// (18, 25, 'local_g1_2')
// (18, 25, 'lutff_2/in_3')
// (18, 25, 'sp4_h_r_2')
// (19, 25, 'sp4_h_r_15')
// (20, 25, 'sp4_h_r_26')
// (21, 22, 'neigh_op_tnr_5')
// (21, 22, 'sp4_r_v_b_39')
// (21, 23, 'neigh_op_rgt_5')
// (21, 23, 'sp4_r_v_b_26')
// (21, 24, 'neigh_op_bnr_5')
// (21, 24, 'sp4_r_v_b_15')
// (21, 25, 'sp4_h_r_39')
// (21, 25, 'sp4_r_v_b_2')
// (22, 21, 'sp4_v_t_39')
// (22, 22, 'neigh_op_top_5')
// (22, 22, 'sp4_v_b_39')
// (22, 23, 'lutff_5/out')
// (22, 23, 'sp4_v_b_26')
// (22, 24, 'neigh_op_bot_5')
// (22, 24, 'sp4_v_b_15')
// (22, 25, 'sp4_h_l_39')
// (22, 25, 'sp4_v_b_2')
// (23, 22, 'neigh_op_tnl_5')
// (23, 23, 'neigh_op_lft_5')
// (23, 24, 'neigh_op_bnl_5')

reg n1419 = 0;
// (18, 25, 'local_g1_3')
// (18, 25, 'lutff_3/in_3')
// (18, 25, 'sp4_h_r_11')
// (19, 25, 'sp4_h_r_22')
// (20, 25, 'sp4_h_r_35')
// (21, 22, 'neigh_op_tnr_7')
// (21, 22, 'sp4_r_v_b_43')
// (21, 23, 'neigh_op_rgt_7')
// (21, 23, 'sp4_r_v_b_30')
// (21, 24, 'neigh_op_bnr_7')
// (21, 24, 'sp4_r_v_b_19')
// (21, 25, 'sp4_h_r_46')
// (21, 25, 'sp4_r_v_b_6')
// (22, 21, 'sp4_v_t_43')
// (22, 22, 'neigh_op_top_7')
// (22, 22, 'sp4_v_b_43')
// (22, 23, 'lutff_7/out')
// (22, 23, 'sp4_v_b_30')
// (22, 24, 'neigh_op_bot_7')
// (22, 24, 'sp4_v_b_19')
// (22, 25, 'sp4_h_l_46')
// (22, 25, 'sp4_v_b_6')
// (23, 22, 'neigh_op_tnl_7')
// (23, 23, 'neigh_op_lft_7')
// (23, 24, 'neigh_op_bnl_7')

reg n1420 = 0;
// (18, 25, 'local_g1_6')
// (18, 25, 'lutff_3/in_0')
// (18, 25, 'sp4_h_r_6')
// (19, 24, 'neigh_op_tnr_7')
// (19, 25, 'neigh_op_rgt_7')
// (19, 25, 'sp4_h_r_19')
// (19, 26, 'neigh_op_bnr_7')
// (20, 24, 'neigh_op_top_7')
// (20, 25, 'lutff_7/out')
// (20, 25, 'sp4_h_r_30')
// (20, 26, 'neigh_op_bot_7')
// (21, 24, 'neigh_op_tnl_7')
// (21, 25, 'neigh_op_lft_7')
// (21, 25, 'sp4_h_r_43')
// (21, 26, 'neigh_op_bnl_7')
// (22, 25, 'sp4_h_l_43')

reg n1421 = 0;
// (18, 26, 'local_g1_5')
// (18, 26, 'lutff_5/in_3')
// (18, 26, 'sp4_h_r_5')
// (19, 26, 'sp4_h_r_16')
// (20, 26, 'sp4_h_r_29')
// (21, 22, 'neigh_op_tnr_4')
// (21, 23, 'neigh_op_rgt_4')
// (21, 23, 'sp4_r_v_b_40')
// (21, 24, 'neigh_op_bnr_4')
// (21, 24, 'sp4_r_v_b_29')
// (21, 25, 'sp4_r_v_b_16')
// (21, 26, 'sp4_h_r_40')
// (21, 26, 'sp4_r_v_b_5')
// (22, 22, 'neigh_op_top_4')
// (22, 22, 'sp4_v_t_40')
// (22, 23, 'lutff_4/out')
// (22, 23, 'sp4_v_b_40')
// (22, 24, 'neigh_op_bot_4')
// (22, 24, 'sp4_v_b_29')
// (22, 25, 'sp4_v_b_16')
// (22, 26, 'sp4_h_l_40')
// (22, 26, 'sp4_v_b_5')
// (23, 22, 'neigh_op_tnl_4')
// (23, 23, 'neigh_op_lft_4')
// (23, 24, 'neigh_op_bnl_4')

reg n1422 = 0;
// (19, 2, 'sp12_v_t_22')
// (19, 3, 'sp12_v_b_22')
// (19, 4, 'sp12_v_b_21')
// (19, 5, 'sp12_v_b_18')
// (19, 6, 'sp12_v_b_17')
// (19, 7, 'sp12_v_b_14')
// (19, 8, 'sp12_v_b_13')
// (19, 9, 'sp12_v_b_10')
// (19, 10, 'sp12_v_b_9')
// (19, 11, 'sp12_v_b_6')
// (19, 12, 'sp12_v_b_5')
// (19, 13, 'local_g3_2')
// (19, 13, 'lutff_1/in_0')
// (19, 13, 'sp12_v_b_2')
// (19, 14, 'sp12_h_r_1')
// (19, 14, 'sp12_v_b_1')
// (20, 14, 'sp12_h_r_2')
// (21, 14, 'sp12_h_r_5')
// (22, 14, 'sp12_h_r_6')
// (23, 13, 'neigh_op_tnr_1')
// (23, 14, 'neigh_op_rgt_1')
// (23, 14, 'sp12_h_r_9')
// (23, 15, 'neigh_op_bnr_1')
// (24, 13, 'neigh_op_top_1')
// (24, 14, 'lutff_1/out')
// (24, 14, 'sp12_h_r_10')
// (24, 15, 'neigh_op_bot_1')
// (25, 13, 'neigh_op_tnl_1')
// (25, 14, 'neigh_op_lft_1')
// (25, 14, 'sp12_h_r_13')
// (25, 15, 'neigh_op_bnl_1')
// (26, 14, 'sp12_h_r_14')
// (27, 14, 'sp12_h_r_17')
// (28, 14, 'sp12_h_r_18')
// (29, 14, 'sp12_h_r_21')
// (30, 14, 'sp12_h_r_22')
// (31, 14, 'sp12_h_l_22')

reg n1423 = 0;
// (19, 7, 'neigh_op_tnr_6')
// (19, 8, 'local_g2_6')
// (19, 8, 'lutff_3/in_3')
// (19, 8, 'neigh_op_rgt_6')
// (19, 9, 'neigh_op_bnr_6')
// (20, 7, 'neigh_op_top_6')
// (20, 8, 'lutff_6/out')
// (20, 9, 'neigh_op_bot_6')
// (21, 7, 'neigh_op_tnl_6')
// (21, 8, 'neigh_op_lft_6')
// (21, 9, 'neigh_op_bnl_6')

wire n1424;
// (19, 8, 'neigh_op_tnr_7')
// (19, 9, 'neigh_op_rgt_7')
// (19, 10, 'neigh_op_bnr_7')
// (20, 8, 'neigh_op_top_7')
// (20, 9, 'lutff_7/out')
// (20, 10, 'neigh_op_bot_7')
// (21, 8, 'neigh_op_tnl_7')
// (21, 9, 'neigh_op_lft_7')
// (21, 10, 'local_g3_7')
// (21, 10, 'lutff_1/in_3')
// (21, 10, 'neigh_op_bnl_7')

reg n1425 = 0;
// (19, 9, 'neigh_op_tnr_3')
// (19, 10, 'neigh_op_rgt_3')
// (19, 10, 'sp4_h_r_11')
// (19, 11, 'neigh_op_bnr_3')
// (20, 9, 'local_g1_3')
// (20, 9, 'lutff_7/in_3')
// (20, 9, 'neigh_op_top_3')
// (20, 10, 'local_g1_3')
// (20, 10, 'lutff_3/in_3')
// (20, 10, 'lutff_3/out')
// (20, 10, 'sp4_h_r_22')
// (20, 11, 'neigh_op_bot_3')
// (21, 9, 'neigh_op_tnl_3')
// (21, 10, 'local_g2_3')
// (21, 10, 'local_g3_3')
// (21, 10, 'lutff_2/in_1')
// (21, 10, 'lutff_5/in_3')
// (21, 10, 'lutff_7/in_2')
// (21, 10, 'neigh_op_lft_3')
// (21, 10, 'sp4_h_r_35')
// (21, 11, 'neigh_op_bnl_3')
// (22, 10, 'local_g3_6')
// (22, 10, 'lutff_0/in_1')
// (22, 10, 'sp4_h_r_46')
// (23, 10, 'sp4_h_l_46')

reg n1426 = 0;
// (19, 9, 'sp4_r_v_b_46')
// (19, 10, 'neigh_op_tnr_3')
// (19, 10, 'sp4_r_v_b_35')
// (19, 11, 'neigh_op_rgt_3')
// (19, 11, 'sp4_r_v_b_22')
// (19, 12, 'neigh_op_bnr_3')
// (19, 12, 'sp4_r_v_b_11')
// (19, 13, 'sp4_r_v_b_46')
// (19, 14, 'sp4_r_v_b_35')
// (19, 15, 'sp4_r_v_b_22')
// (19, 16, 'sp4_r_v_b_11')
// (20, 8, 'sp4_v_t_46')
// (20, 9, 'sp4_v_b_46')
// (20, 10, 'neigh_op_top_3')
// (20, 10, 'sp4_v_b_35')
// (20, 11, 'lutff_3/out')
// (20, 11, 'sp4_v_b_22')
// (20, 12, 'neigh_op_bot_3')
// (20, 12, 'sp4_v_b_11')
// (20, 12, 'sp4_v_t_46')
// (20, 13, 'sp4_v_b_46')
// (20, 14, 'sp4_v_b_35')
// (20, 15, 'sp4_v_b_22')
// (20, 16, 'sp4_h_r_11')
// (20, 16, 'sp4_v_b_11')
// (21, 10, 'neigh_op_tnl_3')
// (21, 11, 'neigh_op_lft_3')
// (21, 12, 'neigh_op_bnl_3')
// (21, 16, 'sp4_h_r_22')
// (22, 16, 'local_g3_3')
// (22, 16, 'lutff_5/in_1')
// (22, 16, 'sp4_h_r_35')
// (23, 16, 'sp4_h_r_46')
// (24, 16, 'sp4_h_l_46')

reg n1427 = 0;
// (19, 10, 'neigh_op_tnr_0')
// (19, 10, 'sp4_r_v_b_45')
// (19, 11, 'neigh_op_rgt_0')
// (19, 11, 'sp4_r_v_b_32')
// (19, 12, 'neigh_op_bnr_0')
// (19, 12, 'sp4_r_v_b_21')
// (19, 13, 'local_g2_0')
// (19, 13, 'lutff_1/in_3')
// (19, 13, 'sp4_r_v_b_8')
// (20, 9, 'sp4_v_t_45')
// (20, 10, 'neigh_op_top_0')
// (20, 10, 'sp4_v_b_45')
// (20, 11, 'lutff_0/out')
// (20, 11, 'sp4_v_b_32')
// (20, 12, 'neigh_op_bot_0')
// (20, 12, 'sp4_v_b_21')
// (20, 13, 'sp4_v_b_8')
// (21, 10, 'neigh_op_tnl_0')
// (21, 11, 'neigh_op_lft_0')
// (21, 12, 'neigh_op_bnl_0')

reg n1428 = 0;
// (19, 10, 'neigh_op_tnr_1')
// (19, 11, 'neigh_op_rgt_1')
// (19, 12, 'neigh_op_bnr_1')
// (20, 10, 'neigh_op_top_1')
// (20, 10, 'sp4_r_v_b_46')
// (20, 11, 'lutff_1/out')
// (20, 11, 'sp4_r_v_b_35')
// (20, 12, 'neigh_op_bot_1')
// (20, 12, 'sp4_r_v_b_22')
// (20, 13, 'sp4_r_v_b_11')
// (21, 9, 'sp4_v_t_46')
// (21, 10, 'neigh_op_tnl_1')
// (21, 10, 'sp4_v_b_46')
// (21, 11, 'neigh_op_lft_1')
// (21, 11, 'sp4_v_b_35')
// (21, 12, 'neigh_op_bnl_1')
// (21, 12, 'sp4_v_b_22')
// (21, 13, 'local_g1_3')
// (21, 13, 'lutff_5/in_1')
// (21, 13, 'sp4_v_b_11')

reg n1429 = 0;
// (19, 10, 'neigh_op_tnr_2')
// (19, 11, 'neigh_op_rgt_2')
// (19, 12, 'neigh_op_bnr_2')
// (20, 10, 'neigh_op_top_2')
// (20, 11, 'lutff_2/out')
// (20, 11, 'sp4_r_v_b_37')
// (20, 12, 'neigh_op_bot_2')
// (20, 12, 'sp4_r_v_b_24')
// (20, 13, 'sp4_r_v_b_13')
// (20, 14, 'sp4_r_v_b_0')
// (20, 15, 'sp4_r_v_b_45')
// (20, 16, 'sp4_r_v_b_32')
// (20, 17, 'sp4_r_v_b_21')
// (20, 18, 'sp4_r_v_b_8')
// (21, 10, 'neigh_op_tnl_2')
// (21, 10, 'sp4_v_t_37')
// (21, 11, 'neigh_op_lft_2')
// (21, 11, 'sp4_v_b_37')
// (21, 12, 'neigh_op_bnl_2')
// (21, 12, 'sp4_v_b_24')
// (21, 13, 'sp4_v_b_13')
// (21, 14, 'sp4_v_b_0')
// (21, 14, 'sp4_v_t_45')
// (21, 15, 'sp4_v_b_45')
// (21, 16, 'local_g2_0')
// (21, 16, 'lutff_3/in_1')
// (21, 16, 'sp4_v_b_32')
// (21, 17, 'sp4_v_b_21')
// (21, 18, 'sp4_v_b_8')

reg n1430 = 0;
// (19, 10, 'neigh_op_tnr_4')
// (19, 11, 'neigh_op_rgt_4')
// (19, 11, 'sp4_r_v_b_40')
// (19, 12, 'neigh_op_bnr_4')
// (19, 12, 'sp4_r_v_b_29')
// (19, 13, 'sp4_r_v_b_16')
// (19, 14, 'sp4_r_v_b_5')
// (19, 15, 'sp4_r_v_b_36')
// (19, 16, 'sp4_r_v_b_25')
// (19, 17, 'sp4_r_v_b_12')
// (19, 18, 'local_g1_1')
// (19, 18, 'lutff_3/in_1')
// (19, 18, 'sp4_r_v_b_1')
// (20, 10, 'neigh_op_top_4')
// (20, 10, 'sp4_v_t_40')
// (20, 11, 'lutff_4/out')
// (20, 11, 'sp4_v_b_40')
// (20, 12, 'neigh_op_bot_4')
// (20, 12, 'sp4_v_b_29')
// (20, 13, 'sp4_v_b_16')
// (20, 14, 'sp4_v_b_5')
// (20, 14, 'sp4_v_t_36')
// (20, 15, 'sp4_v_b_36')
// (20, 16, 'sp4_v_b_25')
// (20, 17, 'sp4_v_b_12')
// (20, 18, 'sp4_v_b_1')
// (21, 10, 'neigh_op_tnl_4')
// (21, 11, 'neigh_op_lft_4')
// (21, 12, 'neigh_op_bnl_4')

reg n1431 = 0;
// (19, 11, 'neigh_op_tnr_0')
// (19, 12, 'neigh_op_rgt_0')
// (19, 13, 'neigh_op_bnr_0')
// (20, 11, 'neigh_op_top_0')
// (20, 11, 'sp4_r_v_b_44')
// (20, 12, 'lutff_0/out')
// (20, 12, 'sp4_r_v_b_33')
// (20, 13, 'neigh_op_bot_0')
// (20, 13, 'sp4_r_v_b_20')
// (20, 14, 'sp4_r_v_b_9')
// (21, 10, 'sp4_v_t_44')
// (21, 11, 'neigh_op_tnl_0')
// (21, 11, 'sp4_v_b_44')
// (21, 12, 'neigh_op_lft_0')
// (21, 12, 'sp4_v_b_33')
// (21, 13, 'neigh_op_bnl_0')
// (21, 13, 'sp4_v_b_20')
// (21, 14, 'local_g1_1')
// (21, 14, 'lutff_1/in_3')
// (21, 14, 'sp4_v_b_9')

reg n1432 = 0;
// (19, 11, 'neigh_op_tnr_1')
// (19, 12, 'neigh_op_rgt_1')
// (19, 13, 'neigh_op_bnr_1')
// (20, 11, 'neigh_op_top_1')
// (20, 11, 'sp4_r_v_b_46')
// (20, 12, 'lutff_1/out')
// (20, 12, 'sp4_r_v_b_35')
// (20, 13, 'neigh_op_bot_1')
// (20, 13, 'sp4_r_v_b_22')
// (20, 14, 'sp4_r_v_b_11')
// (21, 10, 'sp4_v_t_46')
// (21, 11, 'neigh_op_tnl_1')
// (21, 11, 'sp4_v_b_46')
// (21, 12, 'neigh_op_lft_1')
// (21, 12, 'sp4_v_b_35')
// (21, 13, 'neigh_op_bnl_1')
// (21, 13, 'sp4_v_b_22')
// (21, 14, 'local_g0_3')
// (21, 14, 'lutff_4/in_3')
// (21, 14, 'sp4_v_b_11')

reg n1433 = 0;
// (19, 11, 'neigh_op_tnr_3')
// (19, 12, 'neigh_op_rgt_3')
// (19, 12, 'sp4_h_r_11')
// (19, 13, 'neigh_op_bnr_3')
// (20, 11, 'neigh_op_top_3')
// (20, 12, 'lutff_3/out')
// (20, 12, 'sp4_h_r_22')
// (20, 13, 'neigh_op_bot_3')
// (21, 11, 'neigh_op_tnl_3')
// (21, 12, 'neigh_op_lft_3')
// (21, 12, 'sp4_h_r_35')
// (21, 13, 'neigh_op_bnl_3')
// (22, 12, 'sp4_h_r_46')
// (22, 13, 'local_g3_6')
// (22, 13, 'lutff_1/in_0')
// (22, 13, 'sp4_r_v_b_46')
// (22, 14, 'sp4_r_v_b_35')
// (22, 15, 'sp4_r_v_b_22')
// (22, 16, 'sp4_r_v_b_11')
// (23, 12, 'sp4_h_l_46')
// (23, 12, 'sp4_v_t_46')
// (23, 13, 'sp4_v_b_46')
// (23, 14, 'sp4_v_b_35')
// (23, 15, 'sp4_v_b_22')
// (23, 16, 'sp4_v_b_11')

reg n1434 = 0;
// (19, 11, 'sp4_r_v_b_36')
// (19, 12, 'sp4_r_v_b_25')
// (19, 13, 'local_g2_4')
// (19, 13, 'lutff_5/in_3')
// (19, 13, 'sp4_r_v_b_12')
// (19, 14, 'sp4_r_v_b_1')
// (20, 10, 'sp4_v_t_36')
// (20, 11, 'sp4_v_b_36')
// (20, 12, 'sp4_v_b_25')
// (20, 13, 'sp4_v_b_12')
// (20, 14, 'sp4_h_r_8')
// (20, 14, 'sp4_v_b_1')
// (21, 13, 'neigh_op_tnr_0')
// (21, 14, 'neigh_op_rgt_0')
// (21, 14, 'sp4_h_r_21')
// (21, 15, 'neigh_op_bnr_0')
// (22, 13, 'neigh_op_top_0')
// (22, 14, 'lutff_0/out')
// (22, 14, 'sp4_h_r_32')
// (22, 15, 'neigh_op_bot_0')
// (23, 13, 'neigh_op_tnl_0')
// (23, 14, 'neigh_op_lft_0')
// (23, 14, 'sp4_h_r_45')
// (23, 15, 'neigh_op_bnl_0')
// (24, 14, 'sp4_h_l_45')

wire n1435;
// (19, 12, 'lutff_6/lout')
// (19, 12, 'lutff_7/in_2')

wire n1436;
// (19, 12, 'neigh_op_tnr_0')
// (19, 13, 'neigh_op_rgt_0')
// (19, 14, 'neigh_op_bnr_0')
// (20, 12, 'neigh_op_top_0')
// (20, 13, 'local_g1_0')
// (20, 13, 'lutff_0/out')
// (20, 13, 'lutff_2/in_3')
// (20, 14, 'neigh_op_bot_0')
// (21, 12, 'neigh_op_tnl_0')
// (21, 13, 'neigh_op_lft_0')
// (21, 14, 'neigh_op_bnl_0')

wire n1437;
// (19, 12, 'neigh_op_tnr_2')
// (19, 13, 'local_g1_1')
// (19, 13, 'lutff_3/in_1')
// (19, 13, 'neigh_op_rgt_2')
// (19, 13, 'sp4_h_r_9')
// (19, 14, 'neigh_op_bnr_2')
// (20, 12, 'neigh_op_top_2')
// (20, 13, 'lutff_2/out')
// (20, 13, 'sp4_h_r_20')
// (20, 14, 'neigh_op_bot_2')
// (21, 12, 'neigh_op_tnl_2')
// (21, 13, 'neigh_op_lft_2')
// (21, 13, 'sp4_h_r_33')
// (21, 14, 'neigh_op_bnl_2')
// (22, 13, 'sp4_h_r_44')
// (23, 13, 'sp4_h_l_44')

wire n1438;
// (19, 12, 'neigh_op_tnr_4')
// (19, 13, 'neigh_op_rgt_4')
// (19, 14, 'neigh_op_bnr_4')
// (20, 12, 'neigh_op_top_4')
// (20, 13, 'lutff_4/out')
// (20, 14, 'neigh_op_bot_4')
// (21, 12, 'neigh_op_tnl_4')
// (21, 13, 'local_g0_4')
// (21, 13, 'lutff_3/in_1')
// (21, 13, 'neigh_op_lft_4')
// (21, 14, 'neigh_op_bnl_4')

reg n1439 = 0;
// (19, 12, 'neigh_op_tnr_5')
// (19, 13, 'neigh_op_rgt_5')
// (19, 14, 'neigh_op_bnr_5')
// (20, 12, 'neigh_op_top_5')
// (20, 13, 'local_g1_5')
// (20, 13, 'lutff_1/in_3')
// (20, 13, 'lutff_5/out')
// (20, 14, 'neigh_op_bot_5')
// (21, 12, 'neigh_op_tnl_5')
// (21, 13, 'neigh_op_lft_5')
// (21, 14, 'neigh_op_bnl_5')

wire n1440;
// (19, 12, 'neigh_op_tnr_6')
// (19, 13, 'neigh_op_rgt_6')
// (19, 14, 'neigh_op_bnr_6')
// (20, 12, 'neigh_op_top_6')
// (20, 13, 'local_g3_6')
// (20, 13, 'lutff_4/in_3')
// (20, 13, 'lutff_6/out')
// (20, 14, 'neigh_op_bot_6')
// (21, 12, 'neigh_op_tnl_6')
// (21, 13, 'neigh_op_lft_6')
// (21, 14, 'neigh_op_bnl_6')

reg n1441 = 0;
// (19, 12, 'neigh_op_tnr_7')
// (19, 13, 'neigh_op_rgt_7')
// (19, 14, 'neigh_op_bnr_7')
// (20, 12, 'neigh_op_top_7')
// (20, 13, 'local_g1_7')
// (20, 13, 'lutff_3/in_3')
// (20, 13, 'lutff_7/out')
// (20, 14, 'neigh_op_bot_7')
// (21, 12, 'neigh_op_tnl_7')
// (21, 13, 'neigh_op_lft_7')
// (21, 14, 'neigh_op_bnl_7')

reg n1442 = 0;
// (19, 13, 'local_g2_5')
// (19, 13, 'lutff_6/in_1')
// (19, 13, 'sp4_r_v_b_37')
// (19, 14, 'sp4_r_v_b_24')
// (19, 15, 'neigh_op_tnr_0')
// (19, 15, 'sp4_r_v_b_13')
// (19, 16, 'neigh_op_rgt_0')
// (19, 16, 'sp4_r_v_b_0')
// (19, 17, 'neigh_op_bnr_0')
// (20, 12, 'sp4_v_t_37')
// (20, 13, 'sp4_v_b_37')
// (20, 14, 'sp4_v_b_24')
// (20, 15, 'neigh_op_top_0')
// (20, 15, 'sp4_v_b_13')
// (20, 16, 'lutff_0/out')
// (20, 16, 'sp4_v_b_0')
// (20, 17, 'neigh_op_bot_0')
// (21, 15, 'neigh_op_tnl_0')
// (21, 16, 'neigh_op_lft_0')
// (21, 17, 'neigh_op_bnl_0')

wire n1443;
// (19, 13, 'lutff_1/lout')
// (19, 13, 'lutff_2/in_2')

wire n1444;
// (19, 13, 'lutff_2/lout')
// (19, 13, 'lutff_3/in_2')

wire n1445;
// (19, 13, 'lutff_5/lout')
// (19, 13, 'lutff_6/in_2')

wire n1446;
// (19, 13, 'neigh_op_tnr_5')
// (19, 14, 'neigh_op_rgt_5')
// (19, 15, 'neigh_op_bnr_5')
// (20, 13, 'neigh_op_top_5')
// (20, 14, 'local_g1_5')
// (20, 14, 'lutff_1/in_3')
// (20, 14, 'lutff_5/out')
// (20, 15, 'neigh_op_bot_5')
// (21, 13, 'neigh_op_tnl_5')
// (21, 14, 'neigh_op_lft_5')
// (21, 15, 'neigh_op_bnl_5')

wire n1447;
// (19, 13, 'neigh_op_tnr_6')
// (19, 14, 'neigh_op_rgt_6')
// (19, 15, 'neigh_op_bnr_6')
// (20, 13, 'neigh_op_top_6')
// (20, 14, 'local_g3_6')
// (20, 14, 'lutff_0/in_3')
// (20, 14, 'lutff_6/out')
// (20, 15, 'neigh_op_bot_6')
// (21, 13, 'neigh_op_tnl_6')
// (21, 14, 'neigh_op_lft_6')
// (21, 15, 'neigh_op_bnl_6')

reg n1448 = 0;
// (19, 13, 'sp4_r_v_b_47')
// (19, 14, 'local_g0_1')
// (19, 14, 'lutff_2/in_1')
// (19, 14, 'sp4_r_v_b_34')
// (19, 15, 'neigh_op_tnr_5')
// (19, 15, 'sp4_r_v_b_23')
// (19, 16, 'neigh_op_rgt_5')
// (19, 16, 'sp4_r_v_b_10')
// (19, 17, 'neigh_op_bnr_5')
// (20, 12, 'sp4_v_t_47')
// (20, 13, 'sp4_v_b_47')
// (20, 14, 'sp4_v_b_34')
// (20, 15, 'neigh_op_top_5')
// (20, 15, 'sp4_v_b_23')
// (20, 16, 'lutff_5/out')
// (20, 16, 'sp4_v_b_10')
// (20, 17, 'neigh_op_bot_5')
// (21, 15, 'neigh_op_tnl_5')
// (21, 16, 'neigh_op_lft_5')
// (21, 17, 'neigh_op_bnl_5')

reg n1449 = 0;
// (19, 14, 'local_g1_7')
// (19, 14, 'lutff_1/in_3')
// (19, 14, 'sp4_h_r_7')
// (20, 14, 'sp4_h_r_18')
// (21, 13, 'neigh_op_tnr_5')
// (21, 14, 'neigh_op_rgt_5')
// (21, 14, 'sp4_h_r_31')
// (21, 15, 'neigh_op_bnr_5')
// (22, 13, 'neigh_op_top_5')
// (22, 14, 'lutff_5/out')
// (22, 14, 'sp4_h_r_42')
// (22, 15, 'neigh_op_bot_5')
// (23, 13, 'neigh_op_tnl_5')
// (23, 14, 'neigh_op_lft_5')
// (23, 14, 'sp4_h_l_42')
// (23, 15, 'neigh_op_bnl_5')

wire n1450;
// (19, 14, 'lutff_1/lout')
// (19, 14, 'lutff_2/in_2')

wire n1451;
// (19, 14, 'lutff_3/lout')
// (19, 14, 'lutff_4/in_2')

wire n1452;
// (19, 14, 'lutff_4/lout')
// (19, 14, 'lutff_5/in_2')

wire n1453;
// (19, 14, 'neigh_op_tnr_0')
// (19, 15, 'neigh_op_rgt_0')
// (19, 16, 'neigh_op_bnr_0')
// (19, 18, 'sp4_r_v_b_39')
// (19, 19, 'sp4_r_v_b_26')
// (19, 20, 'sp4_r_v_b_15')
// (19, 21, 'sp4_r_v_b_2')
// (19, 22, 'sp4_r_v_b_39')
// (19, 23, 'sp4_r_v_b_26')
// (19, 24, 'sp4_r_v_b_15')
// (19, 25, 'sp4_r_v_b_2')
// (20, 11, 'sp12_v_t_23')
// (20, 12, 'sp12_v_b_23')
// (20, 13, 'sp12_v_b_20')
// (20, 14, 'neigh_op_top_0')
// (20, 14, 'sp12_v_b_19')
// (20, 15, 'lutff_0/out')
// (20, 15, 'sp12_v_b_16')
// (20, 16, 'neigh_op_bot_0')
// (20, 16, 'sp12_v_b_15')
// (20, 17, 'sp12_v_b_12')
// (20, 17, 'sp4_v_t_39')
// (20, 18, 'sp12_v_b_11')
// (20, 18, 'sp4_v_b_39')
// (20, 19, 'sp12_v_b_8')
// (20, 19, 'sp4_v_b_26')
// (20, 20, 'sp12_v_b_7')
// (20, 20, 'sp4_v_b_15')
// (20, 21, 'sp12_v_b_4')
// (20, 21, 'sp4_v_b_2')
// (20, 21, 'sp4_v_t_39')
// (20, 22, 'sp12_v_b_3')
// (20, 22, 'sp4_v_b_39')
// (20, 23, 'sp12_h_r_0')
// (20, 23, 'sp12_v_b_0')
// (20, 23, 'sp12_v_t_23')
// (20, 23, 'sp4_v_b_26')
// (20, 24, 'sp12_v_b_23')
// (20, 24, 'sp4_v_b_15')
// (20, 25, 'local_g0_2')
// (20, 25, 'lutff_global/cen')
// (20, 25, 'sp12_v_b_20')
// (20, 25, 'sp4_v_b_2')
// (20, 26, 'local_g3_3')
// (20, 26, 'lutff_global/cen')
// (20, 26, 'sp12_v_b_19')
// (20, 27, 'sp12_v_b_16')
// (20, 28, 'sp12_v_b_15')
// (20, 29, 'sp12_v_b_12')
// (20, 30, 'sp12_v_b_11')
// (20, 31, 'sp12_v_b_8')
// (20, 32, 'sp12_v_b_7')
// (20, 33, 'span12_vert_4')
// (21, 14, 'neigh_op_tnl_0')
// (21, 15, 'neigh_op_lft_0')
// (21, 16, 'neigh_op_bnl_0')
// (21, 23, 'local_g1_3')
// (21, 23, 'lutff_global/cen')
// (21, 23, 'sp12_h_r_3')
// (22, 23, 'sp12_h_r_4')
// (23, 23, 'sp12_h_r_7')
// (24, 23, 'sp12_h_r_8')
// (25, 23, 'sp12_h_r_11')
// (26, 23, 'sp12_h_r_12')
// (27, 23, 'sp12_h_r_15')
// (28, 23, 'sp12_h_r_16')
// (29, 23, 'sp12_h_r_19')
// (30, 23, 'sp12_h_r_20')
// (31, 23, 'sp12_h_r_23')
// (32, 23, 'sp12_h_l_23')

wire n1454;
// (19, 14, 'neigh_op_tnr_1')
// (19, 15, 'neigh_op_rgt_1')
// (19, 16, 'neigh_op_bnr_1')
// (20, 14, 'neigh_op_top_1')
// (20, 15, 'lutff_1/out')
// (20, 15, 'sp4_h_r_2')
// (20, 16, 'neigh_op_bot_1')
// (21, 14, 'neigh_op_tnl_1')
// (21, 15, 'neigh_op_lft_1')
// (21, 15, 'sp4_h_r_15')
// (21, 16, 'neigh_op_bnl_1')
// (22, 15, 'sp4_h_r_26')
// (23, 15, 'sp4_h_r_39')
// (23, 16, 'sp4_r_v_b_39')
// (23, 17, 'sp4_r_v_b_26')
// (23, 18, 'sp4_r_v_b_15')
// (23, 19, 'sp4_r_v_b_2')
// (24, 15, 'sp4_h_l_39')
// (24, 15, 'sp4_v_t_39')
// (24, 16, 'sp4_v_b_39')
// (24, 17, 'local_g2_2')
// (24, 17, 'lutff_global/cen')
// (24, 17, 'sp4_v_b_26')
// (24, 18, 'sp4_v_b_15')
// (24, 19, 'sp4_v_b_2')

wire n1455;
// (19, 14, 'neigh_op_tnr_2')
// (19, 15, 'neigh_op_rgt_2')
// (19, 16, 'neigh_op_bnr_2')
// (20, 14, 'neigh_op_top_2')
// (20, 15, 'lutff_2/out')
// (20, 16, 'local_g0_2')
// (20, 16, 'lutff_global/cen')
// (20, 16, 'neigh_op_bot_2')
// (21, 14, 'neigh_op_tnl_2')
// (21, 15, 'neigh_op_lft_2')
// (21, 16, 'neigh_op_bnl_2')

wire n1456;
// (19, 14, 'sp4_r_v_b_37')
// (19, 15, 'sp4_r_v_b_24')
// (19, 16, 'sp4_r_v_b_13')
// (19, 17, 'local_g1_0')
// (19, 17, 'lutff_0/in_1')
// (19, 17, 'sp4_r_v_b_0')
// (20, 13, 'sp4_h_r_6')
// (20, 13, 'sp4_v_t_37')
// (20, 14, 'sp4_v_b_37')
// (20, 15, 'sp4_v_b_24')
// (20, 16, 'sp4_v_b_13')
// (20, 17, 'sp4_v_b_0')
// (21, 12, 'neigh_op_tnr_7')
// (21, 13, 'neigh_op_rgt_7')
// (21, 13, 'sp4_h_r_19')
// (21, 14, 'neigh_op_bnr_7')
// (22, 12, 'neigh_op_top_7')
// (22, 13, 'lutff_7/out')
// (22, 13, 'sp4_h_r_30')
// (22, 14, 'neigh_op_bot_7')
// (23, 12, 'neigh_op_tnl_7')
// (23, 13, 'neigh_op_lft_7')
// (23, 13, 'sp4_h_r_43')
// (23, 14, 'neigh_op_bnl_7')
// (24, 13, 'sp4_h_l_43')

wire n1457;
// (19, 14, 'sp4_r_v_b_41')
// (19, 15, 'sp4_r_v_b_28')
// (19, 16, 'neigh_op_tnr_2')
// (19, 16, 'sp4_r_v_b_17')
// (19, 17, 'neigh_op_rgt_2')
// (19, 17, 'sp4_r_v_b_4')
// (19, 18, 'neigh_op_bnr_2')
// (20, 13, 'sp4_v_t_41')
// (20, 14, 'local_g3_1')
// (20, 14, 'lutff_3/in_1')
// (20, 14, 'sp4_v_b_41')
// (20, 15, 'sp4_v_b_28')
// (20, 16, 'neigh_op_top_2')
// (20, 16, 'sp4_v_b_17')
// (20, 17, 'lutff_2/out')
// (20, 17, 'sp4_v_b_4')
// (20, 18, 'neigh_op_bot_2')
// (21, 16, 'neigh_op_tnl_2')
// (21, 17, 'neigh_op_lft_2')
// (21, 18, 'neigh_op_bnl_2')

reg n1458 = 0;
// (19, 14, 'sp4_r_v_b_42')
// (19, 15, 'neigh_op_tnr_1')
// (19, 15, 'sp4_r_v_b_31')
// (19, 16, 'neigh_op_rgt_1')
// (19, 16, 'sp4_r_v_b_18')
// (19, 17, 'neigh_op_bnr_1')
// (19, 17, 'sp4_r_v_b_7')
// (20, 13, 'sp4_h_r_0')
// (20, 13, 'sp4_v_t_42')
// (20, 14, 'sp4_v_b_42')
// (20, 15, 'neigh_op_top_1')
// (20, 15, 'sp4_v_b_31')
// (20, 16, 'lutff_1/out')
// (20, 16, 'sp4_v_b_18')
// (20, 17, 'neigh_op_bot_1')
// (20, 17, 'sp4_v_b_7')
// (21, 13, 'local_g1_5')
// (21, 13, 'lutff_0/in_0')
// (21, 13, 'sp4_h_r_13')
// (21, 15, 'neigh_op_tnl_1')
// (21, 16, 'neigh_op_lft_1')
// (21, 17, 'neigh_op_bnl_1')
// (22, 13, 'sp4_h_r_24')
// (23, 13, 'sp4_h_r_37')
// (24, 13, 'sp4_h_l_37')

reg n1459 = 0;
// (19, 15, 'local_g0_0')
// (19, 15, 'lutff_1/in_1')
// (19, 15, 'sp12_h_r_0')
// (20, 15, 'sp12_h_r_3')
// (21, 15, 'sp12_h_r_4')
// (22, 14, 'neigh_op_tnr_0')
// (22, 15, 'neigh_op_rgt_0')
// (22, 15, 'sp12_h_r_7')
// (22, 16, 'neigh_op_bnr_0')
// (23, 14, 'neigh_op_top_0')
// (23, 15, 'lutff_0/out')
// (23, 15, 'sp12_h_r_8')
// (23, 16, 'neigh_op_bot_0')
// (24, 14, 'neigh_op_tnl_0')
// (24, 15, 'neigh_op_lft_0')
// (24, 15, 'sp12_h_r_11')
// (24, 16, 'neigh_op_bnl_0')
// (25, 15, 'sp12_h_r_12')
// (26, 15, 'sp12_h_r_15')
// (27, 15, 'sp12_h_r_16')
// (28, 15, 'sp12_h_r_19')
// (29, 15, 'sp12_h_r_20')
// (30, 15, 'sp12_h_r_23')
// (31, 15, 'sp12_h_l_23')

reg n1460 = 0;
// (19, 15, 'local_g1_2')
// (19, 15, 'lutff_6/in_1')
// (19, 15, 'sp4_h_r_2')
// (20, 15, 'sp4_h_r_15')
// (21, 15, 'sp4_h_r_26')
// (22, 12, 'sp4_r_v_b_44')
// (22, 13, 'neigh_op_tnr_2')
// (22, 13, 'sp4_r_v_b_33')
// (22, 14, 'neigh_op_rgt_2')
// (22, 14, 'sp4_r_v_b_20')
// (22, 15, 'neigh_op_bnr_2')
// (22, 15, 'sp4_h_r_39')
// (22, 15, 'sp4_r_v_b_9')
// (23, 11, 'sp4_v_t_44')
// (23, 12, 'sp4_v_b_44')
// (23, 13, 'neigh_op_top_2')
// (23, 13, 'sp4_v_b_33')
// (23, 14, 'lutff_2/out')
// (23, 14, 'sp4_v_b_20')
// (23, 15, 'neigh_op_bot_2')
// (23, 15, 'sp4_h_l_39')
// (23, 15, 'sp4_v_b_9')
// (24, 13, 'neigh_op_tnl_2')
// (24, 14, 'neigh_op_lft_2')
// (24, 15, 'neigh_op_bnl_2')

reg n1461 = 0;
// (19, 15, 'local_g1_5')
// (19, 15, 'lutff_1/in_3')
// (19, 15, 'sp4_h_r_5')
// (20, 15, 'sp4_h_r_16')
// (21, 15, 'sp4_h_r_29')
// (22, 12, 'sp4_r_v_b_40')
// (22, 13, 'neigh_op_tnr_0')
// (22, 13, 'sp4_r_v_b_29')
// (22, 14, 'neigh_op_rgt_0')
// (22, 14, 'sp4_r_v_b_16')
// (22, 15, 'neigh_op_bnr_0')
// (22, 15, 'sp4_h_r_40')
// (22, 15, 'sp4_r_v_b_5')
// (23, 11, 'sp4_v_t_40')
// (23, 12, 'sp4_v_b_40')
// (23, 13, 'neigh_op_top_0')
// (23, 13, 'sp4_v_b_29')
// (23, 14, 'lutff_0/out')
// (23, 14, 'sp4_v_b_16')
// (23, 15, 'neigh_op_bot_0')
// (23, 15, 'sp4_h_l_40')
// (23, 15, 'sp4_v_b_5')
// (24, 13, 'neigh_op_tnl_0')
// (24, 14, 'neigh_op_lft_0')
// (24, 15, 'neigh_op_bnl_0')

reg n1462 = 0;
// (19, 15, 'local_g1_7')
// (19, 15, 'lutff_3/in_1')
// (19, 15, 'sp4_h_r_7')
// (20, 15, 'sp4_h_r_18')
// (21, 15, 'sp4_h_r_31')
// (22, 12, 'sp4_r_v_b_42')
// (22, 13, 'neigh_op_tnr_1')
// (22, 13, 'sp4_r_v_b_31')
// (22, 14, 'neigh_op_rgt_1')
// (22, 14, 'sp4_r_v_b_18')
// (22, 15, 'neigh_op_bnr_1')
// (22, 15, 'sp4_h_r_42')
// (22, 15, 'sp4_r_v_b_7')
// (23, 11, 'sp4_v_t_42')
// (23, 12, 'sp4_v_b_42')
// (23, 13, 'neigh_op_top_1')
// (23, 13, 'sp4_v_b_31')
// (23, 14, 'lutff_1/out')
// (23, 14, 'sp4_v_b_18')
// (23, 15, 'neigh_op_bot_1')
// (23, 15, 'sp4_h_l_42')
// (23, 15, 'sp4_v_b_7')
// (24, 13, 'neigh_op_tnl_1')
// (24, 14, 'neigh_op_lft_1')
// (24, 15, 'neigh_op_bnl_1')

wire n1463;
// (19, 15, 'lutff_1/lout')
// (19, 15, 'lutff_2/in_2')

wire n1464;
// (19, 15, 'lutff_3/lout')
// (19, 15, 'lutff_4/in_2')

wire n1465;
// (19, 15, 'lutff_6/lout')
// (19, 15, 'lutff_7/in_2')

reg n1466 = 0;
// (19, 15, 'neigh_op_tnr_2')
// (19, 16, 'neigh_op_rgt_2')
// (19, 16, 'sp4_h_r_9')
// (19, 17, 'neigh_op_bnr_2')
// (20, 15, 'neigh_op_top_2')
// (20, 16, 'lutff_2/out')
// (20, 16, 'sp4_h_r_20')
// (20, 17, 'neigh_op_bot_2')
// (21, 15, 'neigh_op_tnl_2')
// (21, 16, 'local_g2_1')
// (21, 16, 'lutff_2/in_1')
// (21, 16, 'neigh_op_lft_2')
// (21, 16, 'sp4_h_r_33')
// (21, 17, 'neigh_op_bnl_2')
// (22, 16, 'sp4_h_r_44')
// (23, 16, 'sp4_h_l_44')

reg n1467 = 0;
// (19, 15, 'neigh_op_tnr_3')
// (19, 16, 'neigh_op_rgt_3')
// (19, 16, 'sp4_h_r_11')
// (19, 17, 'neigh_op_bnr_3')
// (20, 15, 'neigh_op_top_3')
// (20, 16, 'lutff_3/out')
// (20, 16, 'sp4_h_r_22')
// (20, 17, 'neigh_op_bot_3')
// (21, 15, 'neigh_op_tnl_3')
// (21, 16, 'neigh_op_lft_3')
// (21, 16, 'sp4_h_r_35')
// (21, 17, 'neigh_op_bnl_3')
// (22, 16, 'local_g3_6')
// (22, 16, 'lutff_2/in_1')
// (22, 16, 'sp4_h_r_46')
// (23, 16, 'sp4_h_l_46')

reg n1468 = 0;
// (19, 15, 'neigh_op_tnr_4')
// (19, 16, 'neigh_op_rgt_4')
// (19, 16, 'sp4_r_v_b_40')
// (19, 17, 'neigh_op_bnr_4')
// (19, 17, 'sp4_r_v_b_29')
// (19, 18, 'local_g3_0')
// (19, 18, 'lutff_2/in_1')
// (19, 18, 'sp4_r_v_b_16')
// (19, 19, 'sp4_r_v_b_5')
// (20, 15, 'neigh_op_top_4')
// (20, 15, 'sp4_v_t_40')
// (20, 16, 'lutff_4/out')
// (20, 16, 'sp4_v_b_40')
// (20, 17, 'neigh_op_bot_4')
// (20, 17, 'sp4_v_b_29')
// (20, 18, 'sp4_v_b_16')
// (20, 19, 'sp4_v_b_5')
// (21, 15, 'neigh_op_tnl_4')
// (21, 16, 'neigh_op_lft_4')
// (21, 17, 'neigh_op_bnl_4')

reg n1469 = 0;
// (19, 16, 'neigh_op_tnr_1')
// (19, 17, 'neigh_op_rgt_1')
// (19, 18, 'neigh_op_bnr_1')
// (20, 16, 'neigh_op_top_1')
// (20, 17, 'local_g2_1')
// (20, 17, 'lutff_0/in_3')
// (20, 17, 'lutff_1/out')
// (20, 18, 'neigh_op_bot_1')
// (21, 16, 'neigh_op_tnl_1')
// (21, 17, 'neigh_op_lft_1')
// (21, 18, 'neigh_op_bnl_1')

reg n1470 = 0;
// (19, 16, 'neigh_op_tnr_3')
// (19, 17, 'neigh_op_rgt_3')
// (19, 18, 'neigh_op_bnr_3')
// (20, 16, 'neigh_op_top_3')
// (20, 17, 'local_g0_3')
// (20, 17, 'lutff_2/in_3')
// (20, 17, 'lutff_3/out')
// (20, 18, 'neigh_op_bot_3')
// (21, 16, 'neigh_op_tnl_3')
// (21, 17, 'neigh_op_lft_3')
// (21, 18, 'neigh_op_bnl_3')

wire n1471;
// (19, 16, 'neigh_op_tnr_4')
// (19, 17, 'neigh_op_rgt_4')
// (19, 18, 'neigh_op_bnr_4')
// (20, 16, 'neigh_op_top_4')
// (20, 17, 'lutff_4/out')
// (20, 17, 'sp4_r_v_b_41')
// (20, 18, 'neigh_op_bot_4')
// (20, 18, 'sp4_r_v_b_28')
// (20, 19, 'sp4_r_v_b_17')
// (20, 20, 'sp4_r_v_b_4')
// (21, 16, 'neigh_op_tnl_4')
// (21, 16, 'sp4_v_t_41')
// (21, 17, 'neigh_op_lft_4')
// (21, 17, 'sp4_v_b_41')
// (21, 18, 'neigh_op_bnl_4')
// (21, 18, 'sp4_v_b_28')
// (21, 19, 'local_g0_1')
// (21, 19, 'lutff_0/in_1')
// (21, 19, 'sp4_v_b_17')
// (21, 20, 'sp4_v_b_4')

reg n1472 = 0;
// (19, 16, 'neigh_op_tnr_5')
// (19, 17, 'neigh_op_rgt_5')
// (19, 18, 'neigh_op_bnr_5')
// (20, 16, 'neigh_op_top_5')
// (20, 17, 'local_g2_5')
// (20, 17, 'lutff_4/in_3')
// (20, 17, 'lutff_5/out')
// (20, 18, 'neigh_op_bot_5')
// (21, 16, 'neigh_op_tnl_5')
// (21, 17, 'neigh_op_lft_5')
// (21, 18, 'neigh_op_bnl_5')

wire n1473;
// (19, 16, 'neigh_op_tnr_6')
// (19, 17, 'neigh_op_rgt_6')
// (19, 17, 'sp4_h_r_1')
// (19, 18, 'neigh_op_bnr_6')
// (20, 16, 'neigh_op_top_6')
// (20, 17, 'lutff_6/out')
// (20, 17, 'sp4_h_r_12')
// (20, 18, 'neigh_op_bot_6')
// (21, 16, 'neigh_op_tnl_6')
// (21, 17, 'neigh_op_lft_6')
// (21, 17, 'sp4_h_r_25')
// (21, 18, 'neigh_op_bnl_6')
// (22, 17, 'local_g3_4')
// (22, 17, 'lutff_2/in_1')
// (22, 17, 'sp4_h_r_36')
// (23, 17, 'sp4_h_l_36')

reg n1474 = 0;
// (19, 16, 'neigh_op_tnr_7')
// (19, 17, 'neigh_op_rgt_7')
// (19, 18, 'neigh_op_bnr_7')
// (20, 16, 'neigh_op_top_7')
// (20, 17, 'local_g2_7')
// (20, 17, 'lutff_6/in_3')
// (20, 17, 'lutff_7/out')
// (20, 18, 'neigh_op_bot_7')
// (21, 16, 'neigh_op_tnl_7')
// (21, 17, 'neigh_op_lft_7')
// (21, 18, 'neigh_op_bnl_7')

wire n1475;
// (19, 17, 'local_g0_0')
// (19, 17, 'lutff_5/in_1')
// (19, 17, 'sp4_h_r_0')
// (20, 16, 'neigh_op_tnr_4')
// (20, 17, 'neigh_op_rgt_4')
// (20, 17, 'sp4_h_r_13')
// (20, 18, 'neigh_op_bnr_4')
// (21, 16, 'neigh_op_top_4')
// (21, 17, 'lutff_4/out')
// (21, 17, 'sp4_h_r_24')
// (21, 18, 'neigh_op_bot_4')
// (22, 16, 'neigh_op_tnl_4')
// (22, 17, 'neigh_op_lft_4')
// (22, 17, 'sp4_h_r_37')
// (22, 18, 'neigh_op_bnl_4')
// (23, 17, 'sp4_h_l_37')

wire n1476;
// (19, 17, 'lutff_0/lout')
// (19, 17, 'lutff_1/in_2')

wire n1477;
// (19, 17, 'lutff_1/lout')
// (19, 17, 'lutff_2/in_2')

wire n1478;
// (19, 17, 'lutff_4/lout')
// (19, 17, 'lutff_5/in_2')

wire n1479;
// (19, 17, 'lutff_5/lout')
// (19, 17, 'lutff_6/in_2')

reg n1480 = 0;
// (19, 17, 'neigh_op_tnr_1')
// (19, 18, 'neigh_op_rgt_1')
// (19, 19, 'neigh_op_bnr_1')
// (20, 17, 'neigh_op_top_1')
// (20, 18, 'local_g2_1')
// (20, 18, 'lutff_0/in_3')
// (20, 18, 'lutff_1/out')
// (20, 19, 'neigh_op_bot_1')
// (21, 17, 'neigh_op_tnl_1')
// (21, 18, 'neigh_op_lft_1')
// (21, 19, 'neigh_op_bnl_1')

wire n1481;
// (19, 17, 'neigh_op_tnr_5')
// (19, 18, 'neigh_op_rgt_5')
// (19, 19, 'neigh_op_bnr_5')
// (20, 17, 'neigh_op_top_5')
// (20, 18, 'lutff_5/out')
// (20, 19, 'neigh_op_bot_5')
// (21, 17, 'neigh_op_tnl_5')
// (21, 18, 'neigh_op_lft_5')
// (21, 19, 'local_g3_5')
// (21, 19, 'lutff_1/in_1')
// (21, 19, 'neigh_op_bnl_5')

reg n1482 = 0;
// (19, 17, 'neigh_op_tnr_6')
// (19, 18, 'neigh_op_rgt_6')
// (19, 19, 'neigh_op_bnr_6')
// (20, 17, 'neigh_op_top_6')
// (20, 18, 'local_g2_6')
// (20, 18, 'lutff_5/in_3')
// (20, 18, 'lutff_6/out')
// (20, 19, 'neigh_op_bot_6')
// (21, 17, 'neigh_op_tnl_6')
// (21, 18, 'neigh_op_lft_6')
// (21, 19, 'neigh_op_bnl_6')

reg n1483 = 0;
// (19, 17, 'sp12_h_r_1')
// (20, 17, 'local_g1_2')
// (20, 17, 'lutff_2/in_1')
// (20, 17, 'sp12_h_r_2')
// (21, 17, 'sp12_h_r_5')
// (22, 17, 'sp12_h_r_6')
// (23, 16, 'neigh_op_tnr_1')
// (23, 17, 'neigh_op_rgt_1')
// (23, 17, 'sp12_h_r_9')
// (23, 18, 'neigh_op_bnr_1')
// (24, 16, 'neigh_op_top_1')
// (24, 17, 'lutff_1/out')
// (24, 17, 'sp12_h_r_10')
// (24, 18, 'neigh_op_bot_1')
// (25, 16, 'neigh_op_tnl_1')
// (25, 17, 'neigh_op_lft_1')
// (25, 17, 'sp12_h_r_13')
// (25, 18, 'neigh_op_bnl_1')
// (26, 17, 'sp12_h_r_14')
// (27, 17, 'sp12_h_r_17')
// (28, 17, 'sp12_h_r_18')
// (29, 17, 'sp12_h_r_21')
// (30, 17, 'sp12_h_r_22')
// (31, 17, 'sp12_h_l_22')

reg n1484 = 0;
// (19, 17, 'sp4_h_r_4')
// (20, 17, 'sp4_h_r_17')
// (21, 17, 'local_g3_4')
// (21, 17, 'lutff_0/in_1')
// (21, 17, 'sp4_h_r_28')
// (22, 14, 'sp4_r_v_b_46')
// (22, 15, 'neigh_op_tnr_3')
// (22, 15, 'sp4_r_v_b_35')
// (22, 16, 'neigh_op_rgt_3')
// (22, 16, 'sp4_r_v_b_22')
// (22, 17, 'neigh_op_bnr_3')
// (22, 17, 'sp4_h_r_41')
// (22, 17, 'sp4_r_v_b_11')
// (23, 13, 'sp4_v_t_46')
// (23, 14, 'sp4_v_b_46')
// (23, 15, 'neigh_op_top_3')
// (23, 15, 'sp4_v_b_35')
// (23, 16, 'lutff_3/out')
// (23, 16, 'sp4_v_b_22')
// (23, 17, 'neigh_op_bot_3')
// (23, 17, 'sp4_h_l_41')
// (23, 17, 'sp4_v_b_11')
// (24, 15, 'neigh_op_tnl_3')
// (24, 16, 'neigh_op_lft_3')
// (24, 17, 'neigh_op_bnl_3')

reg n1485 = 0;
// (19, 17, 'sp4_h_r_6')
// (20, 17, 'sp4_h_r_19')
// (21, 17, 'local_g3_6')
// (21, 17, 'lutff_6/in_1')
// (21, 17, 'sp4_h_r_30')
// (22, 14, 'sp4_r_v_b_36')
// (22, 15, 'neigh_op_tnr_6')
// (22, 15, 'sp4_r_v_b_25')
// (22, 16, 'neigh_op_rgt_6')
// (22, 16, 'sp4_r_v_b_12')
// (22, 17, 'neigh_op_bnr_6')
// (22, 17, 'sp4_h_r_43')
// (22, 17, 'sp4_r_v_b_1')
// (23, 13, 'sp4_v_t_36')
// (23, 14, 'sp4_v_b_36')
// (23, 15, 'neigh_op_top_6')
// (23, 15, 'sp4_v_b_25')
// (23, 16, 'lutff_6/out')
// (23, 16, 'sp4_v_b_12')
// (23, 17, 'neigh_op_bot_6')
// (23, 17, 'sp4_h_l_43')
// (23, 17, 'sp4_v_b_1')
// (24, 15, 'neigh_op_tnl_6')
// (24, 16, 'neigh_op_lft_6')
// (24, 17, 'neigh_op_bnl_6')

reg n1486 = 0;
// (19, 17, 'sp4_r_v_b_44')
// (19, 18, 'neigh_op_tnr_2')
// (19, 18, 'sp4_r_v_b_33')
// (19, 19, 'neigh_op_rgt_2')
// (19, 19, 'sp4_r_v_b_20')
// (19, 20, 'neigh_op_bnr_2')
// (19, 20, 'sp4_r_v_b_9')
// (20, 16, 'sp4_v_t_44')
// (20, 17, 'sp4_v_b_44')
// (20, 18, 'neigh_op_top_2')
// (20, 18, 'sp4_v_b_33')
// (20, 19, 'lutff_2/out')
// (20, 19, 'sp4_v_b_20')
// (20, 20, 'neigh_op_bot_2')
// (20, 20, 'sp4_h_r_3')
// (20, 20, 'sp4_v_b_9')
// (21, 18, 'neigh_op_tnl_2')
// (21, 19, 'neigh_op_lft_2')
// (21, 20, 'neigh_op_bnl_2')
// (21, 20, 'sp4_h_r_14')
// (22, 20, 'local_g3_3')
// (22, 20, 'lutff_7/in_3')
// (22, 20, 'sp4_h_r_27')
// (23, 20, 'sp4_h_r_38')
// (24, 20, 'sp4_h_l_38')

wire n1487;
// (19, 18, 'lutff_1/lout')
// (19, 18, 'lutff_2/in_2')

wire n1488;
// (19, 18, 'lutff_3/lout')
// (19, 18, 'lutff_4/in_2')

wire n1489;
// (19, 18, 'lutff_4/lout')
// (19, 18, 'lutff_5/in_2')

reg n1490 = 0;
// (19, 18, 'neigh_op_tnr_1')
// (19, 19, 'neigh_op_rgt_1')
// (19, 20, 'neigh_op_bnr_1')
// (20, 18, 'neigh_op_top_1')
// (20, 18, 'sp4_r_v_b_46')
// (20, 19, 'lutff_1/out')
// (20, 19, 'sp4_r_v_b_35')
// (20, 20, 'neigh_op_bot_1')
// (20, 20, 'sp4_r_v_b_22')
// (20, 21, 'sp4_r_v_b_11')
// (21, 17, 'sp4_v_t_46')
// (21, 18, 'neigh_op_tnl_1')
// (21, 18, 'sp4_v_b_46')
// (21, 19, 'neigh_op_lft_1')
// (21, 19, 'sp4_v_b_35')
// (21, 20, 'neigh_op_bnl_1')
// (21, 20, 'sp4_v_b_22')
// (21, 21, 'local_g1_3')
// (21, 21, 'lutff_5/in_3')
// (21, 21, 'sp4_v_b_11')

reg n1491 = 0;
// (19, 18, 'sp4_h_r_5')
// (20, 18, 'sp4_h_r_16')
// (21, 18, 'sp4_h_r_29')
// (22, 11, 'neigh_op_tnr_4')
// (22, 11, 'sp4_r_v_b_37')
// (22, 12, 'neigh_op_rgt_4')
// (22, 12, 'sp4_r_v_b_24')
// (22, 13, 'neigh_op_bnr_4')
// (22, 13, 'sp4_r_v_b_13')
// (22, 14, 'sp4_r_v_b_0')
// (22, 15, 'sp4_r_v_b_37')
// (22, 16, 'sp4_r_v_b_24')
// (22, 17, 'sp4_r_v_b_13')
// (22, 18, 'local_g3_0')
// (22, 18, 'lutff_2/in_1')
// (22, 18, 'sp4_h_r_40')
// (22, 18, 'sp4_r_v_b_0')
// (23, 10, 'sp4_v_t_37')
// (23, 11, 'neigh_op_top_4')
// (23, 11, 'sp4_v_b_37')
// (23, 12, 'lutff_4/out')
// (23, 12, 'sp4_v_b_24')
// (23, 13, 'neigh_op_bot_4')
// (23, 13, 'sp4_v_b_13')
// (23, 14, 'sp4_v_b_0')
// (23, 14, 'sp4_v_t_37')
// (23, 15, 'sp4_v_b_37')
// (23, 16, 'sp4_v_b_24')
// (23, 17, 'sp4_v_b_13')
// (23, 18, 'sp4_h_l_40')
// (23, 18, 'sp4_v_b_0')
// (24, 11, 'neigh_op_tnl_4')
// (24, 12, 'neigh_op_lft_4')
// (24, 13, 'neigh_op_bnl_4')

wire n1492;
// (19, 18, 'sp4_r_v_b_37')
// (19, 19, 'sp4_r_v_b_24')
// (19, 20, 'neigh_op_tnr_0')
// (19, 20, 'sp4_r_v_b_13')
// (19, 21, 'neigh_op_rgt_0')
// (19, 21, 'sp4_r_v_b_0')
// (19, 22, 'neigh_op_bnr_0')
// (20, 17, 'sp4_h_r_5')
// (20, 17, 'sp4_v_t_37')
// (20, 18, 'sp4_v_b_37')
// (20, 19, 'sp4_v_b_24')
// (20, 20, 'neigh_op_top_0')
// (20, 20, 'sp4_v_b_13')
// (20, 21, 'lutff_0/out')
// (20, 21, 'sp4_v_b_0')
// (20, 22, 'neigh_op_bot_0')
// (21, 17, 'sp4_h_r_16')
// (21, 20, 'neigh_op_tnl_0')
// (21, 21, 'neigh_op_lft_0')
// (21, 22, 'neigh_op_bnl_0')
// (22, 17, 'local_g2_5')
// (22, 17, 'lutff_2/in_3')
// (22, 17, 'sp4_h_r_29')
// (23, 17, 'sp4_h_r_40')
// (24, 17, 'sp4_h_l_40')

reg n1493 = 0;
// (19, 19, 'neigh_op_tnr_1')
// (19, 20, 'neigh_op_rgt_1')
// (19, 21, 'neigh_op_bnr_1')
// (20, 19, 'neigh_op_top_1')
// (20, 20, 'lutff_1/out')
// (20, 21, 'neigh_op_bot_1')
// (21, 19, 'neigh_op_tnl_1')
// (21, 20, 'neigh_op_lft_1')
// (21, 21, 'local_g2_1')
// (21, 21, 'lutff_0/in_1')
// (21, 21, 'neigh_op_bnl_1')

wire n1494;
// (19, 19, 'sp12_h_r_0')
// (19, 20, 'sp4_r_v_b_44')
// (19, 21, 'local_g2_1')
// (19, 21, 'lutff_7/in_2')
// (19, 21, 'sp4_r_v_b_33')
// (19, 22, 'sp4_r_v_b_20')
// (19, 23, 'sp4_r_v_b_9')
// (20, 19, 'sp12_h_r_3')
// (20, 19, 'sp4_h_r_3')
// (20, 19, 'sp4_v_t_44')
// (20, 20, 'sp4_v_b_44')
// (20, 21, 'sp4_v_b_33')
// (20, 22, 'sp4_v_b_20')
// (20, 23, 'sp4_v_b_9')
// (21, 19, 'sp12_h_r_4')
// (21, 19, 'sp4_h_r_14')
// (22, 19, 'sp12_h_r_7')
// (22, 19, 'sp4_h_r_27')
// (23, 19, 'sp12_h_r_8')
// (23, 19, 'sp4_h_r_38')
// (24, 19, 'sp12_h_r_11')
// (24, 19, 'sp4_h_l_38')
// (25, 19, 'sp12_h_r_12')
// (26, 19, 'sp12_h_r_15')
// (27, 19, 'sp12_h_r_16')
// (28, 19, 'sp12_h_r_19')
// (29, 19, 'sp12_h_r_20')
// (30, 19, 'sp12_h_r_23')
// (30, 32, 'neigh_op_tnr_2')
// (30, 32, 'neigh_op_tnr_6')
// (31, 19, 'sp12_h_l_23')
// (31, 19, 'sp12_v_t_23')
// (31, 20, 'sp12_v_b_23')
// (31, 21, 'sp12_v_b_20')
// (31, 22, 'sp12_v_b_19')
// (31, 23, 'sp12_v_b_16')
// (31, 24, 'sp12_v_b_15')
// (31, 25, 'sp12_v_b_12')
// (31, 26, 'sp12_v_b_11')
// (31, 27, 'sp12_v_b_8')
// (31, 28, 'sp12_v_b_7')
// (31, 29, 'sp12_v_b_4')
// (31, 30, 'sp12_v_b_3')
// (31, 31, 'sp12_v_b_0')
// (31, 31, 'sp12_v_t_23')
// (31, 32, 'neigh_op_top_2')
// (31, 32, 'neigh_op_top_6')
// (31, 32, 'sp12_v_b_23')
// (31, 33, 'io_1/D_IN_0')
// (31, 33, 'span12_vert_20')
// (32, 32, 'neigh_op_tnl_2')
// (32, 32, 'neigh_op_tnl_6')

wire n1495;
// (19, 19, 'sp4_r_v_b_44')
// (19, 20, 'neigh_op_tnr_2')
// (19, 20, 'sp4_r_v_b_33')
// (19, 21, 'neigh_op_rgt_2')
// (19, 21, 'sp4_r_v_b_20')
// (19, 22, 'neigh_op_bnr_2')
// (19, 22, 'sp4_r_v_b_9')
// (20, 18, 'sp4_h_r_9')
// (20, 18, 'sp4_v_t_44')
// (20, 19, 'sp4_v_b_44')
// (20, 20, 'neigh_op_top_2')
// (20, 20, 'sp4_v_b_33')
// (20, 21, 'lutff_2/out')
// (20, 21, 'sp4_v_b_20')
// (20, 22, 'neigh_op_bot_2')
// (20, 22, 'sp4_v_b_9')
// (21, 18, 'sp4_h_r_20')
// (21, 20, 'neigh_op_tnl_2')
// (21, 21, 'neigh_op_lft_2')
// (21, 22, 'neigh_op_bnl_2')
// (22, 18, 'local_g2_1')
// (22, 18, 'lutff_4/in_3')
// (22, 18, 'sp4_h_r_33')
// (23, 18, 'sp4_h_r_44')
// (24, 18, 'sp4_h_l_44')

reg n1496 = 0;
// (19, 20, 'neigh_op_tnr_1')
// (19, 21, 'neigh_op_rgt_1')
// (19, 22, 'neigh_op_bnr_1')
// (20, 20, 'neigh_op_top_1')
// (20, 21, 'local_g2_1')
// (20, 21, 'lutff_0/in_3')
// (20, 21, 'lutff_1/out')
// (20, 22, 'neigh_op_bot_1')
// (21, 20, 'neigh_op_tnl_1')
// (21, 21, 'neigh_op_lft_1')
// (21, 22, 'neigh_op_bnl_1')

reg n1497 = 0;
// (19, 20, 'neigh_op_tnr_3')
// (19, 21, 'neigh_op_rgt_3')
// (19, 22, 'neigh_op_bnr_3')
// (20, 20, 'neigh_op_top_3')
// (20, 21, 'local_g0_3')
// (20, 21, 'lutff_2/in_3')
// (20, 21, 'lutff_3/out')
// (20, 22, 'neigh_op_bot_3')
// (21, 20, 'neigh_op_tnl_3')
// (21, 21, 'neigh_op_lft_3')
// (21, 22, 'neigh_op_bnl_3')

reg n1498 = 0;
// (19, 20, 'neigh_op_tnr_5')
// (19, 21, 'neigh_op_rgt_5')
// (19, 22, 'neigh_op_bnr_5')
// (20, 20, 'neigh_op_top_5')
// (20, 21, 'local_g2_5')
// (20, 21, 'lutff_4/in_3')
// (20, 21, 'lutff_5/out')
// (20, 22, 'neigh_op_bot_5')
// (21, 20, 'neigh_op_tnl_5')
// (21, 21, 'neigh_op_lft_5')
// (21, 22, 'neigh_op_bnl_5')

reg n1499 = 0;
// (19, 20, 'neigh_op_tnr_7')
// (19, 21, 'neigh_op_rgt_7')
// (19, 22, 'neigh_op_bnr_7')
// (20, 20, 'neigh_op_top_7')
// (20, 21, 'local_g2_7')
// (20, 21, 'lutff_6/in_3')
// (20, 21, 'lutff_7/out')
// (20, 22, 'neigh_op_bot_7')
// (21, 20, 'neigh_op_tnl_7')
// (21, 21, 'neigh_op_lft_7')
// (21, 22, 'neigh_op_bnl_7')

wire n1500;
// (19, 20, 'sp4_r_v_b_36')
// (19, 21, 'local_g1_1')
// (19, 21, 'lutff_1/in_1')
// (19, 21, 'sp4_r_v_b_25')
// (19, 22, 'sp4_r_v_b_12')
// (19, 23, 'sp4_r_v_b_1')
// (20, 19, 'sp4_v_t_36')
// (20, 20, 'sp4_v_b_36')
// (20, 21, 'sp4_v_b_25')
// (20, 22, 'sp4_v_b_12')
// (20, 23, 'sp4_h_r_8')
// (20, 23, 'sp4_v_b_1')
// (21, 23, 'sp4_h_r_21')
// (22, 23, 'sp4_h_r_32')
// (23, 23, 'sp4_h_r_45')
// (24, 23, 'sp4_h_l_45')
// (24, 23, 'sp4_h_r_8')
// (25, 23, 'sp4_h_r_21')
// (26, 23, 'sp4_h_r_32')
// (27, 23, 'sp4_h_r_45')
// (27, 24, 'sp4_r_v_b_45')
// (27, 25, 'sp4_r_v_b_32')
// (27, 26, 'sp4_r_v_b_21')
// (27, 27, 'sp4_r_v_b_8')
// (27, 32, 'neigh_op_tnr_2')
// (27, 32, 'neigh_op_tnr_6')
// (28, 23, 'sp12_v_t_23')
// (28, 23, 'sp4_h_l_45')
// (28, 23, 'sp4_v_t_45')
// (28, 24, 'sp12_v_b_23')
// (28, 24, 'sp4_v_b_45')
// (28, 25, 'sp12_v_b_20')
// (28, 25, 'sp4_v_b_32')
// (28, 26, 'sp12_v_b_19')
// (28, 26, 'sp4_v_b_21')
// (28, 27, 'sp12_v_b_16')
// (28, 27, 'sp4_v_b_8')
// (28, 28, 'sp12_v_b_15')
// (28, 29, 'sp12_v_b_12')
// (28, 30, 'sp12_v_b_11')
// (28, 31, 'sp12_v_b_8')
// (28, 32, 'neigh_op_top_2')
// (28, 32, 'neigh_op_top_6')
// (28, 32, 'sp12_v_b_7')
// (28, 33, 'io_1/D_IN_0')
// (28, 33, 'span12_vert_4')
// (29, 32, 'neigh_op_tnl_2')
// (29, 32, 'neigh_op_tnl_6')

wire n1501;
// (19, 20, 'sp4_r_v_b_37')
// (19, 21, 'sp4_r_v_b_24')
// (19, 22, 'neigh_op_tnr_0')
// (19, 22, 'sp4_r_v_b_13')
// (19, 23, 'neigh_op_rgt_0')
// (19, 23, 'sp4_r_v_b_0')
// (19, 24, 'local_g0_0')
// (19, 24, 'local_g1_0')
// (19, 24, 'lutff_0/in_0')
// (19, 24, 'lutff_1/in_0')
// (19, 24, 'lutff_2/in_0')
// (19, 24, 'lutff_3/in_0')
// (19, 24, 'lutff_4/in_0')
// (19, 24, 'lutff_5/in_0')
// (19, 24, 'lutff_6/in_0')
// (19, 24, 'lutff_7/in_0')
// (19, 24, 'neigh_op_bnr_0')
// (20, 19, 'sp4_v_t_37')
// (20, 20, 'sp4_v_b_37')
// (20, 21, 'sp4_v_b_24')
// (20, 22, 'local_g1_5')
// (20, 22, 'lutff_6/in_2')
// (20, 22, 'neigh_op_top_0')
// (20, 22, 'sp4_v_b_13')
// (20, 23, 'lutff_0/out')
// (20, 23, 'sp4_v_b_0')
// (20, 24, 'neigh_op_bot_0')
// (21, 22, 'neigh_op_tnl_0')
// (21, 23, 'neigh_op_lft_0')
// (21, 24, 'neigh_op_bnl_0')

wire n1502;
// (19, 21, 'local_g1_0')
// (19, 21, 'lutff_6/in_1')
// (19, 21, 'sp12_h_r_0')
// (20, 21, 'sp12_h_r_3')
// (21, 21, 'sp12_h_r_4')
// (22, 21, 'sp12_h_r_7')
// (23, 21, 'sp12_h_r_8')
// (24, 21, 'sp12_h_r_11')
// (25, 21, 'sp12_h_r_12')
// (26, 21, 'sp12_h_r_15')
// (27, 21, 'sp12_h_r_16')
// (28, 21, 'sp12_h_r_19')
// (29, 21, 'sp12_h_r_20')
// (30, 21, 'sp12_h_r_23')
// (30, 32, 'neigh_op_tnr_0')
// (30, 32, 'neigh_op_tnr_4')
// (31, 21, 'sp12_h_l_23')
// (31, 21, 'sp12_v_t_23')
// (31, 22, 'sp12_v_b_23')
// (31, 23, 'sp12_v_b_20')
// (31, 24, 'sp12_v_b_19')
// (31, 25, 'sp12_v_b_16')
// (31, 26, 'sp12_v_b_15')
// (31, 27, 'sp12_v_b_12')
// (31, 28, 'sp12_v_b_11')
// (31, 29, 'sp12_v_b_8')
// (31, 30, 'sp12_v_b_7')
// (31, 31, 'sp12_v_b_4')
// (31, 32, 'neigh_op_top_0')
// (31, 32, 'neigh_op_top_4')
// (31, 32, 'sp12_v_b_3')
// (31, 33, 'io_0/D_IN_0')
// (31, 33, 'span12_vert_0')
// (32, 32, 'neigh_op_tnl_0')
// (32, 32, 'neigh_op_tnl_4')

wire n1503;
// (19, 21, 'neigh_op_tnr_0')
// (19, 22, 'neigh_op_rgt_0')
// (19, 23, 'neigh_op_bnr_0')
// (20, 21, 'neigh_op_top_0')
// (20, 22, 'local_g1_0')
// (20, 22, 'lutff_0/out')
// (20, 22, 'lutff_4/in_3')
// (20, 23, 'neigh_op_bot_0')
// (21, 21, 'neigh_op_tnl_0')
// (21, 22, 'neigh_op_lft_0')
// (21, 23, 'neigh_op_bnl_0')

reg n1504 = 0;
// (19, 21, 'neigh_op_tnr_2')
// (19, 22, 'neigh_op_rgt_2')
// (19, 23, 'neigh_op_bnr_2')
// (20, 21, 'neigh_op_top_2')
// (20, 22, 'local_g2_2')
// (20, 22, 'local_g3_2')
// (20, 22, 'lutff_2/in_0')
// (20, 22, 'lutff_2/out')
// (20, 22, 'lutff_3/in_0')
// (20, 23, 'neigh_op_bot_2')
// (21, 21, 'neigh_op_tnl_2')
// (21, 22, 'neigh_op_lft_2')
// (21, 23, 'neigh_op_bnl_2')

reg n1505 = 0;
// (19, 21, 'sp4_h_r_1')
// (20, 21, 'local_g1_4')
// (20, 21, 'lutff_6/in_1')
// (20, 21, 'sp4_h_r_12')
// (21, 21, 'sp4_h_r_25')
// (22, 18, 'sp4_r_v_b_36')
// (22, 19, 'neigh_op_tnr_6')
// (22, 19, 'sp4_r_v_b_25')
// (22, 20, 'neigh_op_rgt_6')
// (22, 20, 'sp4_r_v_b_12')
// (22, 21, 'neigh_op_bnr_6')
// (22, 21, 'sp4_h_r_36')
// (22, 21, 'sp4_r_v_b_1')
// (23, 17, 'sp4_v_t_36')
// (23, 18, 'sp4_v_b_36')
// (23, 19, 'neigh_op_top_6')
// (23, 19, 'sp4_v_b_25')
// (23, 20, 'lutff_6/out')
// (23, 20, 'sp4_v_b_12')
// (23, 21, 'neigh_op_bot_6')
// (23, 21, 'sp4_h_l_36')
// (23, 21, 'sp4_v_b_1')
// (24, 19, 'neigh_op_tnl_6')
// (24, 20, 'neigh_op_lft_6')
// (24, 21, 'neigh_op_bnl_6')

reg n1506 = 0;
// (19, 21, 'sp4_h_r_4')
// (20, 21, 'local_g0_1')
// (20, 21, 'lutff_0/in_1')
// (20, 21, 'sp4_h_r_17')
// (21, 21, 'sp4_h_r_28')
// (22, 18, 'sp4_r_v_b_46')
// (22, 19, 'neigh_op_tnr_3')
// (22, 19, 'sp4_r_v_b_35')
// (22, 20, 'neigh_op_rgt_3')
// (22, 20, 'sp4_r_v_b_22')
// (22, 21, 'neigh_op_bnr_3')
// (22, 21, 'sp4_h_r_41')
// (22, 21, 'sp4_r_v_b_11')
// (23, 17, 'sp4_v_t_46')
// (23, 18, 'sp4_v_b_46')
// (23, 19, 'neigh_op_top_3')
// (23, 19, 'sp4_v_b_35')
// (23, 20, 'lutff_3/out')
// (23, 20, 'sp4_v_b_22')
// (23, 21, 'neigh_op_bot_3')
// (23, 21, 'sp4_h_l_41')
// (23, 21, 'sp4_v_b_11')
// (24, 19, 'neigh_op_tnl_3')
// (24, 20, 'neigh_op_lft_3')
// (24, 21, 'neigh_op_bnl_3')

reg n1507 = 0;
// (19, 21, 'sp4_r_v_b_40')
// (19, 22, 'sp4_r_v_b_29')
// (19, 23, 'sp4_r_v_b_16')
// (19, 24, 'sp4_r_v_b_5')
// (20, 20, 'sp4_h_r_5')
// (20, 20, 'sp4_v_t_40')
// (20, 21, 'local_g3_0')
// (20, 21, 'lutff_2/in_1')
// (20, 21, 'sp4_v_b_40')
// (20, 22, 'sp4_v_b_29')
// (20, 23, 'sp4_v_b_16')
// (20, 24, 'sp4_v_b_5')
// (21, 20, 'sp4_h_r_16')
// (22, 19, 'neigh_op_tnr_4')
// (22, 20, 'neigh_op_rgt_4')
// (22, 20, 'sp4_h_r_29')
// (22, 21, 'neigh_op_bnr_4')
// (23, 19, 'neigh_op_top_4')
// (23, 20, 'lutff_4/out')
// (23, 20, 'sp4_h_r_40')
// (23, 21, 'neigh_op_bot_4')
// (24, 19, 'neigh_op_tnl_4')
// (24, 20, 'neigh_op_lft_4')
// (24, 20, 'sp4_h_l_40')
// (24, 21, 'neigh_op_bnl_4')

reg n1508 = 0;
// (19, 21, 'sp4_r_v_b_42')
// (19, 22, 'sp4_r_v_b_31')
// (19, 23, 'sp4_r_v_b_18')
// (19, 24, 'sp4_r_v_b_7')
// (20, 20, 'sp4_h_r_7')
// (20, 20, 'sp4_v_t_42')
// (20, 21, 'local_g3_2')
// (20, 21, 'lutff_4/in_1')
// (20, 21, 'sp4_v_b_42')
// (20, 22, 'sp4_v_b_31')
// (20, 23, 'sp4_v_b_18')
// (20, 24, 'sp4_v_b_7')
// (21, 20, 'sp4_h_r_18')
// (22, 19, 'neigh_op_tnr_5')
// (22, 20, 'neigh_op_rgt_5')
// (22, 20, 'sp4_h_r_31')
// (22, 21, 'neigh_op_bnr_5')
// (23, 19, 'neigh_op_top_5')
// (23, 20, 'lutff_5/out')
// (23, 20, 'sp4_h_r_42')
// (23, 21, 'neigh_op_bot_5')
// (24, 19, 'neigh_op_tnl_5')
// (24, 20, 'neigh_op_lft_5')
// (24, 20, 'sp4_h_l_42')
// (24, 21, 'neigh_op_bnl_5')

reg n1509 = 0;
// (19, 21, 'sp4_r_v_b_43')
// (19, 22, 'sp4_r_v_b_30')
// (19, 23, 'sp4_r_v_b_19')
// (19, 24, 'neigh_op_tnr_3')
// (19, 24, 'sp4_r_v_b_6')
// (19, 25, 'neigh_op_rgt_3')
// (19, 25, 'sp4_r_v_b_38')
// (19, 26, 'neigh_op_bnr_3')
// (19, 26, 'sp4_r_v_b_27')
// (19, 27, 'sp4_r_v_b_14')
// (19, 28, 'sp4_r_v_b_3')
// (20, 20, 'sp4_h_r_6')
// (20, 20, 'sp4_v_t_43')
// (20, 21, 'sp4_v_b_43')
// (20, 22, 'sp4_v_b_30')
// (20, 23, 'sp4_v_b_19')
// (20, 24, 'neigh_op_top_3')
// (20, 24, 'sp4_v_b_6')
// (20, 24, 'sp4_v_t_38')
// (20, 25, 'lutff_3/out')
// (20, 25, 'sp4_v_b_38')
// (20, 26, 'neigh_op_bot_3')
// (20, 26, 'sp4_v_b_27')
// (20, 27, 'sp4_v_b_14')
// (20, 28, 'sp4_v_b_3')
// (21, 20, 'sp4_h_r_19')
// (21, 24, 'neigh_op_tnl_3')
// (21, 25, 'neigh_op_lft_3')
// (21, 26, 'neigh_op_bnl_3')
// (22, 20, 'local_g3_6')
// (22, 20, 'lutff_6/in_1')
// (22, 20, 'sp4_h_r_30')
// (23, 20, 'sp4_h_r_43')
// (24, 20, 'sp4_h_l_43')

wire n1510;
// (19, 22, 'carry_in_mux')
// (19, 22, 'lutff_0/in_3')

wire n1511;
// (19, 22, 'lutff_0/cout')
// (19, 22, 'lutff_1/in_3')

wire n1512;
// (19, 22, 'lutff_1/cout')
// (19, 22, 'lutff_2/in_3')

wire n1513;
// (19, 22, 'lutff_2/cout')
// (19, 22, 'lutff_3/in_3')

wire n1514;
// (19, 22, 'lutff_3/cout')
// (19, 22, 'lutff_4/in_3')

wire n1515;
// (19, 22, 'lutff_4/cout')
// (19, 22, 'lutff_5/in_3')

wire n1516;
// (19, 22, 'lutff_5/cout')
// (19, 22, 'lutff_6/in_3')

wire n1517;
// (19, 22, 'lutff_6/cout')
// (19, 22, 'lutff_7/in_3')

reg n1518 = 0;
// (19, 22, 'neigh_op_tnr_2')
// (19, 23, 'neigh_op_rgt_2')
// (19, 23, 'sp4_r_v_b_36')
// (19, 24, 'neigh_op_bnr_2')
// (19, 24, 'sp4_r_v_b_25')
// (19, 25, 'sp4_r_v_b_12')
// (19, 26, 'sp4_r_v_b_1')
// (20, 22, 'neigh_op_top_2')
// (20, 22, 'sp4_v_t_36')
// (20, 23, 'lutff_2/out')
// (20, 23, 'sp4_v_b_36')
// (20, 24, 'local_g2_1')
// (20, 24, 'lutff_1/in_0')
// (20, 24, 'neigh_op_bot_2')
// (20, 24, 'sp4_v_b_25')
// (20, 25, 'sp4_v_b_12')
// (20, 26, 'sp4_v_b_1')
// (21, 22, 'neigh_op_tnl_2')
// (21, 23, 'neigh_op_lft_2')
// (21, 24, 'neigh_op_bnl_2')

reg n1519 = 0;
// (19, 22, 'neigh_op_tnr_3')
// (19, 23, 'neigh_op_rgt_3')
// (19, 24, 'neigh_op_bnr_3')
// (20, 22, 'neigh_op_top_3')
// (20, 23, 'lutff_3/out')
// (20, 24, 'local_g1_3')
// (20, 24, 'lutff_1/in_3')
// (20, 24, 'neigh_op_bot_3')
// (21, 22, 'neigh_op_tnl_3')
// (21, 23, 'neigh_op_lft_3')
// (21, 24, 'neigh_op_bnl_3')

reg n1520 = 0;
// (19, 22, 'neigh_op_tnr_5')
// (19, 23, 'neigh_op_rgt_5')
// (19, 24, 'neigh_op_bnr_5')
// (20, 22, 'neigh_op_top_5')
// (20, 23, 'lutff_5/out')
// (20, 24, 'local_g1_5')
// (20, 24, 'lutff_2/in_0')
// (20, 24, 'neigh_op_bot_5')
// (21, 22, 'neigh_op_tnl_5')
// (21, 23, 'neigh_op_lft_5')
// (21, 24, 'neigh_op_bnl_5')

reg n1521 = 0;
// (19, 22, 'neigh_op_tnr_6')
// (19, 23, 'neigh_op_rgt_6')
// (19, 24, 'neigh_op_bnr_6')
// (20, 22, 'neigh_op_top_6')
// (20, 23, 'lutff_6/out')
// (20, 24, 'local_g0_6')
// (20, 24, 'lutff_2/in_2')
// (20, 24, 'neigh_op_bot_6')
// (21, 22, 'neigh_op_tnl_6')
// (21, 23, 'neigh_op_lft_6')
// (21, 24, 'neigh_op_bnl_6')

wire n1522;
// (19, 23, 'neigh_op_tnr_1')
// (19, 24, 'neigh_op_rgt_1')
// (19, 25, 'neigh_op_bnr_1')
// (20, 23, 'local_g0_1')
// (20, 23, 'lutff_0/in_1')
// (20, 23, 'neigh_op_top_1')
// (20, 24, 'lutff_1/out')
// (20, 25, 'neigh_op_bot_1')
// (21, 23, 'neigh_op_tnl_1')
// (21, 24, 'neigh_op_lft_1')
// (21, 25, 'neigh_op_bnl_1')

wire n1523;
// (19, 23, 'neigh_op_tnr_2')
// (19, 24, 'neigh_op_rgt_2')
// (19, 25, 'neigh_op_bnr_2')
// (20, 23, 'local_g1_2')
// (20, 23, 'lutff_0/in_3')
// (20, 23, 'neigh_op_top_2')
// (20, 24, 'lutff_2/out')
// (20, 25, 'neigh_op_bot_2')
// (21, 23, 'neigh_op_tnl_2')
// (21, 24, 'neigh_op_lft_2')
// (21, 25, 'neigh_op_bnl_2')

wire n1524;
// (19, 23, 'neigh_op_tnr_7')
// (19, 24, 'neigh_op_rgt_7')
// (19, 25, 'neigh_op_bnr_7')
// (20, 23, 'local_g1_7')
// (20, 23, 'lutff_0/in_0')
// (20, 23, 'neigh_op_top_7')
// (20, 24, 'lutff_7/out')
// (20, 25, 'neigh_op_bot_7')
// (21, 23, 'neigh_op_tnl_7')
// (21, 24, 'neigh_op_lft_7')
// (21, 25, 'neigh_op_bnl_7')

wire n1525;
// (19, 24, 'carry_in_mux')
// (19, 24, 'lutff_0/in_3')

wire n1526;
// (19, 24, 'lutff_0/cout')
// (19, 24, 'lutff_1/in_3')

wire n1527;
// (19, 24, 'lutff_1/cout')
// (19, 24, 'lutff_2/in_3')

wire n1528;
// (19, 24, 'lutff_2/cout')
// (19, 24, 'lutff_3/in_3')

wire n1529;
// (19, 24, 'lutff_3/cout')
// (19, 24, 'lutff_4/in_3')

wire n1530;
// (19, 24, 'lutff_4/cout')
// (19, 24, 'lutff_5/in_3')

wire n1531;
// (19, 24, 'lutff_5/cout')
// (19, 24, 'lutff_6/in_3')

wire n1532;
// (19, 24, 'lutff_6/cout')
// (19, 24, 'lutff_7/in_3')

reg n1533 = 0;
// (19, 24, 'neigh_op_tnr_2')
// (19, 25, 'neigh_op_rgt_2')
// (19, 26, 'neigh_op_bnr_2')
// (20, 22, 'sp4_r_v_b_40')
// (20, 23, 'sp4_r_v_b_29')
// (20, 24, 'neigh_op_top_2')
// (20, 24, 'sp4_r_v_b_16')
// (20, 25, 'lutff_2/out')
// (20, 25, 'sp4_r_v_b_5')
// (20, 26, 'neigh_op_bot_2')
// (21, 21, 'sp4_v_t_40')
// (21, 22, 'local_g3_0')
// (21, 22, 'lutff_0/in_1')
// (21, 22, 'sp4_v_b_40')
// (21, 23, 'sp4_v_b_29')
// (21, 24, 'neigh_op_tnl_2')
// (21, 24, 'sp4_v_b_16')
// (21, 25, 'neigh_op_lft_2')
// (21, 25, 'sp4_v_b_5')
// (21, 26, 'neigh_op_bnl_2')

wire n1534;
// (20, 9, 'neigh_op_tnr_0')
// (20, 10, 'neigh_op_rgt_0')
// (20, 11, 'neigh_op_bnr_0')
// (21, 9, 'neigh_op_top_0')
// (21, 10, 'local_g2_0')
// (21, 10, 'lutff_0/out')
// (21, 10, 'lutff_7/in_3')
// (21, 11, 'neigh_op_bot_0')
// (22, 9, 'neigh_op_tnl_0')
// (22, 10, 'neigh_op_lft_0')
// (22, 11, 'neigh_op_bnl_0')

reg n1535 = 0;
// (20, 9, 'neigh_op_tnr_2')
// (20, 10, 'neigh_op_rgt_2')
// (20, 11, 'neigh_op_bnr_2')
// (21, 9, 'neigh_op_top_2')
// (21, 10, 'local_g3_2')
// (21, 10, 'lutff_0/in_1')
// (21, 10, 'lutff_2/in_3')
// (21, 10, 'lutff_2/out')
// (21, 10, 'lutff_4/in_3')
// (21, 11, 'neigh_op_bot_2')
// (22, 9, 'neigh_op_tnl_2')
// (22, 10, 'local_g0_2')
// (22, 10, 'lutff_0/in_2')
// (22, 10, 'neigh_op_lft_2')
// (22, 11, 'neigh_op_bnl_2')

wire n1536;
// (20, 9, 'neigh_op_tnr_3')
// (20, 10, 'neigh_op_rgt_3')
// (20, 11, 'neigh_op_bnr_3')
// (21, 9, 'neigh_op_top_3')
// (21, 10, 'local_g0_3')
// (21, 10, 'lutff_0/in_3')
// (21, 10, 'lutff_3/out')
// (21, 10, 'lutff_5/in_0')
// (21, 11, 'neigh_op_bot_3')
// (22, 9, 'neigh_op_tnl_3')
// (22, 10, 'neigh_op_lft_3')
// (22, 11, 'neigh_op_bnl_3')

wire n1537;
// (20, 9, 'neigh_op_tnr_5')
// (20, 10, 'local_g2_5')
// (20, 10, 'lutff_0/in_1')
// (20, 10, 'neigh_op_rgt_5')
// (20, 11, 'neigh_op_bnr_5')
// (21, 9, 'neigh_op_top_5')
// (21, 10, 'lutff_5/out')
// (21, 11, 'neigh_op_bot_5')
// (22, 9, 'neigh_op_tnl_5')
// (22, 10, 'local_g0_5')
// (22, 10, 'lutff_7/in_0')
// (22, 10, 'neigh_op_lft_5')
// (22, 11, 'neigh_op_bnl_5')

reg n1538 = 0;
// (20, 9, 'neigh_op_tnr_6')
// (20, 10, 'neigh_op_rgt_6')
// (20, 11, 'neigh_op_bnr_6')
// (21, 9, 'neigh_op_top_6')
// (21, 10, 'local_g2_6')
// (21, 10, 'lutff_3/in_1')
// (21, 10, 'lutff_6/in_0')
// (21, 10, 'lutff_6/out')
// (21, 11, 'neigh_op_bot_6')
// (22, 9, 'neigh_op_tnl_6')
// (22, 10, 'local_g0_6')
// (22, 10, 'lutff_5/in_1')
// (22, 10, 'neigh_op_lft_6')
// (22, 11, 'neigh_op_bnl_6')

wire n1539;
// (20, 9, 'neigh_op_tnr_7')
// (20, 10, 'local_g2_7')
// (20, 10, 'lutff_0/in_3')
// (20, 10, 'neigh_op_rgt_7')
// (20, 11, 'neigh_op_bnr_7')
// (21, 9, 'neigh_op_top_7')
// (21, 10, 'lutff_7/out')
// (21, 11, 'neigh_op_bot_7')
// (22, 9, 'neigh_op_tnl_7')
// (22, 10, 'neigh_op_lft_7')
// (22, 11, 'neigh_op_bnl_7')

reg n1540 = 0;
// (20, 10, 'local_g0_6')
// (20, 10, 'lutff_0/in_0')
// (20, 10, 'sp4_h_r_6')
// (21, 9, 'neigh_op_tnr_7')
// (21, 10, 'local_g2_7')
// (21, 10, 'lutff_1/in_0')
// (21, 10, 'lutff_6/in_1')
// (21, 10, 'neigh_op_rgt_7')
// (21, 10, 'sp4_h_r_19')
// (21, 11, 'neigh_op_bnr_7')
// (22, 9, 'neigh_op_top_7')
// (22, 10, 'local_g3_7')
// (22, 10, 'lutff_7/in_1')
// (22, 10, 'lutff_7/out')
// (22, 10, 'sp4_h_r_30')
// (22, 11, 'neigh_op_bot_7')
// (23, 9, 'neigh_op_tnl_7')
// (23, 10, 'neigh_op_lft_7')
// (23, 10, 'sp4_h_r_43')
// (23, 11, 'neigh_op_bnl_7')
// (24, 10, 'sp4_h_l_43')

reg n1541 = 0;
// (20, 10, 'neigh_op_tnr_1')
// (20, 10, 'sp4_r_v_b_47')
// (20, 11, 'neigh_op_rgt_1')
// (20, 11, 'sp4_r_v_b_34')
// (20, 12, 'neigh_op_bnr_1')
// (20, 12, 'sp4_r_v_b_23')
// (20, 13, 'local_g2_2')
// (20, 13, 'lutff_1/in_1')
// (20, 13, 'sp4_r_v_b_10')
// (21, 9, 'sp4_v_t_47')
// (21, 10, 'neigh_op_top_1')
// (21, 10, 'sp4_v_b_47')
// (21, 11, 'lutff_1/out')
// (21, 11, 'sp4_v_b_34')
// (21, 12, 'neigh_op_bot_1')
// (21, 12, 'sp4_v_b_23')
// (21, 13, 'sp4_v_b_10')
// (22, 10, 'neigh_op_tnl_1')
// (22, 11, 'neigh_op_lft_1')
// (22, 12, 'neigh_op_bnl_1')

reg n1542 = 0;
// (20, 10, 'neigh_op_tnr_2')
// (20, 11, 'neigh_op_rgt_2')
// (20, 11, 'sp4_r_v_b_36')
// (20, 12, 'neigh_op_bnr_2')
// (20, 12, 'sp4_r_v_b_25')
// (20, 13, 'local_g2_4')
// (20, 13, 'lutff_3/in_1')
// (20, 13, 'sp4_r_v_b_12')
// (20, 14, 'sp4_r_v_b_1')
// (21, 10, 'neigh_op_top_2')
// (21, 10, 'sp4_v_t_36')
// (21, 11, 'lutff_2/out')
// (21, 11, 'sp4_v_b_36')
// (21, 12, 'neigh_op_bot_2')
// (21, 12, 'sp4_v_b_25')
// (21, 13, 'sp4_v_b_12')
// (21, 14, 'sp4_v_b_1')
// (22, 10, 'neigh_op_tnl_2')
// (22, 11, 'neigh_op_lft_2')
// (22, 12, 'neigh_op_bnl_2')

reg n1543 = 0;
// (20, 10, 'neigh_op_tnr_3')
// (20, 11, 'neigh_op_rgt_3')
// (20, 12, 'neigh_op_bnr_3')
// (21, 10, 'neigh_op_top_3')
// (21, 10, 'sp12_v_t_22')
// (21, 11, 'lutff_3/out')
// (21, 11, 'sp12_v_b_22')
// (21, 12, 'neigh_op_bot_3')
// (21, 12, 'sp12_v_b_21')
// (21, 13, 'sp12_v_b_18')
// (21, 14, 'sp12_v_b_17')
// (21, 15, 'local_g2_6')
// (21, 15, 'lutff_1/in_1')
// (21, 15, 'sp12_v_b_14')
// (21, 16, 'sp12_v_b_13')
// (21, 17, 'sp12_v_b_10')
// (21, 18, 'sp12_v_b_9')
// (21, 19, 'sp12_v_b_6')
// (21, 20, 'sp12_v_b_5')
// (21, 21, 'sp12_v_b_2')
// (21, 22, 'sp12_v_b_1')
// (22, 10, 'neigh_op_tnl_3')
// (22, 11, 'neigh_op_lft_3')
// (22, 12, 'neigh_op_bnl_3')

reg n1544 = 0;
// (20, 10, 'neigh_op_tnr_4')
// (20, 11, 'neigh_op_rgt_4')
// (20, 12, 'neigh_op_bnr_4')
// (21, 3, 'sp12_v_t_23')
// (21, 4, 'sp12_v_b_23')
// (21, 5, 'sp12_v_b_20')
// (21, 6, 'sp12_v_b_19')
// (21, 7, 'sp12_v_b_16')
// (21, 8, 'sp12_v_b_15')
// (21, 9, 'sp12_v_b_12')
// (21, 10, 'neigh_op_top_4')
// (21, 10, 'sp12_v_b_11')
// (21, 11, 'lutff_4/out')
// (21, 11, 'sp12_v_b_8')
// (21, 12, 'neigh_op_bot_4')
// (21, 12, 'sp12_v_b_7')
// (21, 13, 'sp12_v_b_4')
// (21, 14, 'sp12_v_b_3')
// (21, 15, 'local_g2_0')
// (21, 15, 'lutff_3/in_1')
// (21, 15, 'sp12_v_b_0')
// (22, 10, 'neigh_op_tnl_4')
// (22, 11, 'neigh_op_lft_4')
// (22, 12, 'neigh_op_bnl_4')

reg n1545 = 0;
// (20, 11, 'neigh_op_tnr_0')
// (20, 11, 'sp4_r_v_b_45')
// (20, 12, 'neigh_op_rgt_0')
// (20, 12, 'sp4_r_v_b_32')
// (20, 13, 'neigh_op_bnr_0')
// (20, 13, 'sp4_r_v_b_21')
// (20, 14, 'sp4_r_v_b_8')
// (21, 10, 'sp4_v_t_45')
// (21, 11, 'neigh_op_top_0')
// (21, 11, 'sp4_v_b_45')
// (21, 12, 'lutff_0/out')
// (21, 12, 'sp4_v_b_32')
// (21, 13, 'neigh_op_bot_0')
// (21, 13, 'sp4_v_b_21')
// (21, 14, 'local_g0_0')
// (21, 14, 'lutff_1/in_1')
// (21, 14, 'sp4_v_b_8')
// (22, 11, 'neigh_op_tnl_0')
// (22, 12, 'neigh_op_lft_0')
// (22, 13, 'neigh_op_bnl_0')

reg n1546 = 0;
// (20, 11, 'neigh_op_tnr_1')
// (20, 12, 'neigh_op_rgt_1')
// (20, 13, 'neigh_op_bnr_1')
// (21, 11, 'neigh_op_top_1')
// (21, 11, 'sp4_r_v_b_46')
// (21, 12, 'lutff_1/out')
// (21, 12, 'sp4_r_v_b_35')
// (21, 13, 'neigh_op_bot_1')
// (21, 13, 'sp4_r_v_b_22')
// (21, 14, 'local_g2_3')
// (21, 14, 'lutff_4/in_1')
// (21, 14, 'sp4_r_v_b_11')
// (22, 10, 'sp4_v_t_46')
// (22, 11, 'neigh_op_tnl_1')
// (22, 11, 'sp4_v_b_46')
// (22, 12, 'neigh_op_lft_1')
// (22, 12, 'sp4_v_b_35')
// (22, 13, 'neigh_op_bnl_1')
// (22, 13, 'sp4_v_b_22')
// (22, 14, 'sp4_v_b_11')

reg n1547 = 0;
// (20, 11, 'neigh_op_tnr_2')
// (20, 12, 'neigh_op_rgt_2')
// (20, 12, 'sp4_r_v_b_36')
// (20, 13, 'neigh_op_bnr_2')
// (20, 13, 'sp4_r_v_b_25')
// (20, 14, 'sp4_r_v_b_12')
// (20, 15, 'sp4_r_v_b_1')
// (21, 11, 'neigh_op_top_2')
// (21, 11, 'sp4_v_t_36')
// (21, 12, 'lutff_2/out')
// (21, 12, 'sp4_v_b_36')
// (21, 13, 'neigh_op_bot_2')
// (21, 13, 'sp4_v_b_25')
// (21, 14, 'local_g0_4')
// (21, 14, 'lutff_7/in_1')
// (21, 14, 'sp4_v_b_12')
// (21, 15, 'sp4_v_b_1')
// (22, 11, 'neigh_op_tnl_2')
// (22, 12, 'neigh_op_lft_2')
// (22, 13, 'neigh_op_bnl_2')

reg n1548 = 0;
// (20, 11, 'neigh_op_tnr_3')
// (20, 12, 'neigh_op_rgt_3')
// (20, 13, 'neigh_op_bnr_3')
// (21, 11, 'neigh_op_top_3')
// (21, 12, 'lutff_3/out')
// (21, 13, 'neigh_op_bot_3')
// (22, 11, 'neigh_op_tnl_3')
// (22, 12, 'neigh_op_lft_3')
// (22, 13, 'local_g3_3')
// (22, 13, 'lutff_1/in_3')
// (22, 13, 'neigh_op_bnl_3')

reg n1549 = 0;
// (20, 11, 'neigh_op_tnr_4')
// (20, 12, 'neigh_op_rgt_4')
// (20, 13, 'neigh_op_bnr_4')
// (21, 11, 'neigh_op_top_4')
// (21, 12, 'lutff_4/out')
// (21, 13, 'neigh_op_bot_4')
// (22, 11, 'neigh_op_tnl_4')
// (22, 12, 'neigh_op_lft_4')
// (22, 13, 'local_g3_4')
// (22, 13, 'lutff_4/in_1')
// (22, 13, 'neigh_op_bnl_4')

reg n1550 = 0;
// (20, 11, 'neigh_op_tnr_5')
// (20, 12, 'neigh_op_rgt_5')
// (20, 13, 'neigh_op_bnr_5')
// (21, 11, 'neigh_op_top_5')
// (21, 12, 'lutff_5/out')
// (21, 13, 'neigh_op_bot_5')
// (22, 11, 'neigh_op_tnl_5')
// (22, 12, 'neigh_op_lft_5')
// (22, 13, 'local_g3_5')
// (22, 13, 'lutff_7/in_1')
// (22, 13, 'neigh_op_bnl_5')

wire n1551;
// (20, 12, 'neigh_op_tnr_0')
// (20, 13, 'neigh_op_rgt_0')
// (20, 14, 'local_g1_0')
// (20, 14, 'lutff_6/in_3')
// (20, 14, 'neigh_op_bnr_0')
// (21, 12, 'neigh_op_top_0')
// (21, 13, 'lutff_0/out')
// (21, 14, 'neigh_op_bot_0')
// (22, 12, 'neigh_op_tnl_0')
// (22, 13, 'neigh_op_lft_0')
// (22, 14, 'neigh_op_bnl_0')

wire n1552;
// (20, 12, 'neigh_op_tnr_3')
// (20, 13, 'neigh_op_rgt_3')
// (20, 14, 'neigh_op_bnr_3')
// (21, 12, 'neigh_op_top_3')
// (21, 12, 'sp12_v_t_22')
// (21, 13, 'lutff_3/out')
// (21, 13, 'sp12_v_b_22')
// (21, 14, 'neigh_op_bot_3')
// (21, 14, 'sp12_v_b_21')
// (21, 15, 'sp12_v_b_18')
// (21, 16, 'sp12_v_b_17')
// (21, 17, 'sp12_v_b_14')
// (21, 18, 'sp12_v_b_13')
// (21, 19, 'local_g2_2')
// (21, 19, 'lutff_5/in_1')
// (21, 19, 'sp12_v_b_10')
// (21, 20, 'sp12_v_b_9')
// (21, 21, 'sp12_v_b_6')
// (21, 22, 'sp12_v_b_5')
// (21, 23, 'sp12_v_b_2')
// (21, 24, 'sp12_v_b_1')
// (22, 12, 'neigh_op_tnl_3')
// (22, 13, 'neigh_op_lft_3')
// (22, 14, 'neigh_op_bnl_3')

reg n1553 = 0;
// (20, 12, 'neigh_op_tnr_4')
// (20, 13, 'neigh_op_rgt_4')
// (20, 14, 'neigh_op_bnr_4')
// (21, 12, 'neigh_op_top_4')
// (21, 13, 'local_g1_4')
// (21, 13, 'lutff_0/in_1')
// (21, 13, 'lutff_4/out')
// (21, 14, 'neigh_op_bot_4')
// (22, 12, 'neigh_op_tnl_4')
// (22, 13, 'neigh_op_lft_4')
// (22, 14, 'neigh_op_bnl_4')

wire n1554;
// (20, 12, 'neigh_op_tnr_6')
// (20, 13, 'neigh_op_rgt_6')
// (20, 14, 'neigh_op_bnr_6')
// (21, 12, 'neigh_op_top_6')
// (21, 13, 'local_g2_6')
// (21, 13, 'lutff_3/in_3')
// (21, 13, 'lutff_6/out')
// (21, 14, 'neigh_op_bot_6')
// (22, 12, 'neigh_op_tnl_6')
// (22, 13, 'neigh_op_lft_6')
// (22, 14, 'neigh_op_bnl_6')

wire n1555;
// (20, 12, 'neigh_op_tnr_7')
// (20, 13, 'neigh_op_rgt_7')
// (20, 14, 'neigh_op_bnr_7')
// (21, 12, 'neigh_op_top_7')
// (21, 13, 'local_g2_7')
// (21, 13, 'lutff_0/in_3')
// (21, 13, 'lutff_7/out')
// (21, 14, 'neigh_op_bot_7')
// (22, 12, 'neigh_op_tnl_7')
// (22, 13, 'neigh_op_lft_7')
// (22, 14, 'neigh_op_bnl_7')

reg n1556 = 0;
// (20, 12, 'sp4_r_v_b_47')
// (20, 13, 'sp4_r_v_b_34')
// (20, 14, 'sp4_r_v_b_23')
// (20, 15, 'sp4_r_v_b_10')
// (21, 11, 'sp4_h_r_10')
// (21, 11, 'sp4_v_t_47')
// (21, 12, 'sp4_v_b_47')
// (21, 13, 'sp4_v_b_34')
// (21, 14, 'sp4_v_b_23')
// (21, 15, 'local_g1_2')
// (21, 15, 'lutff_6/in_1')
// (21, 15, 'sp4_v_b_10')
// (22, 10, 'neigh_op_tnr_1')
// (22, 11, 'neigh_op_rgt_1')
// (22, 11, 'sp4_h_r_23')
// (22, 12, 'neigh_op_bnr_1')
// (23, 10, 'neigh_op_top_1')
// (23, 11, 'lutff_1/out')
// (23, 11, 'sp4_h_r_34')
// (23, 12, 'neigh_op_bot_1')
// (24, 10, 'neigh_op_tnl_1')
// (24, 11, 'neigh_op_lft_1')
// (24, 11, 'sp4_h_r_47')
// (24, 12, 'neigh_op_bnl_1')
// (25, 11, 'sp4_h_l_47')

wire n1557;
// (20, 13, 'lutff_1/lout')
// (20, 13, 'lutff_2/in_2')

wire n1558;
// (20, 13, 'lutff_3/lout')
// (20, 13, 'lutff_4/in_2')

reg n1559 = 0;
// (20, 13, 'neigh_op_tnr_2')
// (20, 14, 'neigh_op_rgt_2')
// (20, 15, 'neigh_op_bnr_2')
// (21, 13, 'neigh_op_top_2')
// (21, 14, 'local_g3_2')
// (21, 14, 'lutff_0/in_3')
// (21, 14, 'lutff_2/out')
// (21, 15, 'neigh_op_bot_2')
// (22, 13, 'neigh_op_tnl_2')
// (22, 14, 'neigh_op_lft_2')
// (22, 15, 'neigh_op_bnl_2')

wire n1560;
// (20, 13, 'neigh_op_tnr_4')
// (20, 14, 'local_g2_4')
// (20, 14, 'lutff_0/in_0')
// (20, 14, 'neigh_op_rgt_4')
// (20, 15, 'neigh_op_bnr_4')
// (21, 13, 'neigh_op_top_4')
// (21, 14, 'lutff_4/out')
// (21, 15, 'neigh_op_bot_4')
// (22, 13, 'neigh_op_tnl_4')
// (22, 14, 'neigh_op_lft_4')
// (22, 15, 'neigh_op_bnl_4')

reg n1561 = 0;
// (20, 13, 'neigh_op_tnr_5')
// (20, 14, 'neigh_op_rgt_5')
// (20, 15, 'neigh_op_bnr_5')
// (21, 13, 'neigh_op_top_5')
// (21, 14, 'local_g1_5')
// (21, 14, 'lutff_3/in_3')
// (21, 14, 'lutff_5/out')
// (21, 15, 'neigh_op_bot_5')
// (22, 13, 'neigh_op_tnl_5')
// (22, 14, 'neigh_op_lft_5')
// (22, 15, 'neigh_op_bnl_5')

wire n1562;
// (20, 13, 'neigh_op_tnr_7')
// (20, 14, 'neigh_op_rgt_7')
// (20, 15, 'neigh_op_bnr_7')
// (21, 9, 'sp12_v_t_22')
// (21, 10, 'sp12_v_b_22')
// (21, 11, 'sp12_v_b_21')
// (21, 12, 'sp12_v_b_18')
// (21, 13, 'neigh_op_top_7')
// (21, 13, 'sp12_v_b_17')
// (21, 14, 'lutff_7/out')
// (21, 14, 'sp12_v_b_14')
// (21, 15, 'neigh_op_bot_7')
// (21, 15, 'sp12_v_b_13')
// (21, 16, 'sp12_v_b_10')
// (21, 17, 'sp12_v_b_9')
// (21, 18, 'sp12_v_b_6')
// (21, 19, 'local_g2_5')
// (21, 19, 'lutff_4/in_3')
// (21, 19, 'sp12_v_b_5')
// (21, 20, 'sp12_v_b_2')
// (21, 21, 'sp12_v_b_1')
// (22, 13, 'neigh_op_tnl_7')
// (22, 14, 'neigh_op_lft_7')
// (22, 15, 'neigh_op_bnl_7')

reg n1563 = 0;
// (20, 13, 'sp4_h_r_7')
// (21, 13, 'local_g0_2')
// (21, 13, 'lutff_5/in_3')
// (21, 13, 'sp4_h_r_18')
// (22, 13, 'sp4_h_r_31')
// (23, 13, 'neigh_op_tnr_2')
// (23, 13, 'sp4_h_r_42')
// (23, 14, 'neigh_op_rgt_2')
// (23, 14, 'sp4_r_v_b_36')
// (23, 15, 'neigh_op_bnr_2')
// (23, 15, 'sp4_r_v_b_25')
// (23, 16, 'sp4_r_v_b_12')
// (23, 17, 'sp4_r_v_b_1')
// (24, 13, 'neigh_op_top_2')
// (24, 13, 'sp4_h_l_42')
// (24, 13, 'sp4_v_t_36')
// (24, 14, 'lutff_2/out')
// (24, 14, 'sp4_v_b_36')
// (24, 15, 'neigh_op_bot_2')
// (24, 15, 'sp4_v_b_25')
// (24, 16, 'sp4_v_b_12')
// (24, 17, 'sp4_v_b_1')
// (25, 13, 'neigh_op_tnl_2')
// (25, 14, 'neigh_op_lft_2')
// (25, 15, 'neigh_op_bnl_2')

wire n1564;
// (20, 13, 'sp4_r_v_b_45')
// (20, 14, 'local_g0_3')
// (20, 14, 'lutff_4/in_1')
// (20, 14, 'sp4_r_v_b_32')
// (20, 15, 'sp4_r_v_b_21')
// (20, 16, 'sp4_r_v_b_8')
// (20, 21, 'neigh_op_tnr_2')
// (20, 22, 'neigh_op_rgt_2')
// (20, 23, 'neigh_op_bnr_2')
// (21, 12, 'sp12_v_t_23')
// (21, 12, 'sp4_v_t_45')
// (21, 13, 'sp12_v_b_23')
// (21, 13, 'sp4_v_b_45')
// (21, 14, 'sp12_v_b_20')
// (21, 14, 'sp4_v_b_32')
// (21, 15, 'sp12_v_b_19')
// (21, 15, 'sp4_v_b_21')
// (21, 16, 'sp12_v_b_16')
// (21, 16, 'sp4_v_b_8')
// (21, 17, 'sp12_v_b_15')
// (21, 18, 'sp12_v_b_12')
// (21, 19, 'sp12_v_b_11')
// (21, 20, 'sp12_v_b_8')
// (21, 21, 'neigh_op_top_2')
// (21, 21, 'sp12_v_b_7')
// (21, 22, 'lutff_2/out')
// (21, 22, 'sp12_v_b_4')
// (21, 23, 'neigh_op_bot_2')
// (21, 23, 'sp12_v_b_3')
// (21, 24, 'sp12_v_b_0')
// (22, 21, 'neigh_op_tnl_2')
// (22, 22, 'neigh_op_lft_2')
// (22, 23, 'neigh_op_bnl_2')

reg n1565 = 0;
// (20, 14, 'local_g1_4')
// (20, 14, 'lutff_2/in_1')
// (20, 14, 'sp4_h_r_4')
// (21, 14, 'sp4_h_r_17')
// (22, 11, 'neigh_op_tnr_1')
// (22, 12, 'neigh_op_rgt_1')
// (22, 13, 'neigh_op_bnr_1')
// (22, 14, 'sp4_h_r_28')
// (23, 11, 'neigh_op_top_1')
// (23, 11, 'sp4_r_v_b_46')
// (23, 12, 'lutff_1/out')
// (23, 12, 'sp4_r_v_b_35')
// (23, 13, 'neigh_op_bot_1')
// (23, 13, 'sp4_r_v_b_22')
// (23, 14, 'sp4_h_r_41')
// (23, 14, 'sp4_r_v_b_11')
// (24, 10, 'sp4_v_t_46')
// (24, 11, 'neigh_op_tnl_1')
// (24, 11, 'sp4_v_b_46')
// (24, 12, 'neigh_op_lft_1')
// (24, 12, 'sp4_v_b_35')
// (24, 13, 'neigh_op_bnl_1')
// (24, 13, 'sp4_v_b_22')
// (24, 14, 'sp4_h_l_41')
// (24, 14, 'sp4_v_b_11')

wire n1566;
// (20, 14, 'local_g2_5')
// (20, 14, 'lutff_5/in_0')
// (20, 14, 'sp4_r_v_b_37')
// (20, 15, 'sp4_r_v_b_24')
// (20, 16, 'sp4_r_v_b_13')
// (20, 17, 'sp4_r_v_b_0')
// (20, 18, 'sp4_r_v_b_41')
// (20, 19, 'sp4_r_v_b_28')
// (20, 20, 'neigh_op_tnr_2')
// (20, 20, 'sp4_r_v_b_17')
// (20, 21, 'neigh_op_rgt_2')
// (20, 21, 'sp4_r_v_b_4')
// (20, 22, 'neigh_op_bnr_2')
// (21, 13, 'sp4_v_t_37')
// (21, 14, 'sp4_v_b_37')
// (21, 15, 'sp4_v_b_24')
// (21, 16, 'sp4_v_b_13')
// (21, 17, 'sp4_v_b_0')
// (21, 17, 'sp4_v_t_41')
// (21, 18, 'sp4_v_b_41')
// (21, 19, 'sp4_v_b_28')
// (21, 20, 'neigh_op_top_2')
// (21, 20, 'sp4_v_b_17')
// (21, 21, 'lutff_2/out')
// (21, 21, 'sp4_v_b_4')
// (21, 22, 'neigh_op_bot_2')
// (22, 20, 'neigh_op_tnl_2')
// (22, 21, 'neigh_op_lft_2')
// (22, 22, 'neigh_op_bnl_2')

wire n1567;
// (20, 14, 'lutff_0/lout')
// (20, 14, 'lutff_1/in_2')

wire n1568;
// (20, 14, 'lutff_1/lout')
// (20, 14, 'lutff_2/in_2')

wire n1569;
// (20, 14, 'lutff_3/lout')
// (20, 14, 'lutff_4/in_2')

wire n1570;
// (20, 14, 'lutff_4/lout')
// (20, 14, 'lutff_5/in_2')

wire n1571;
// (20, 14, 'neigh_op_tnr_0')
// (20, 15, 'neigh_op_rgt_0')
// (20, 16, 'neigh_op_bnr_0')
// (21, 14, 'neigh_op_top_0')
// (21, 15, 'local_g3_0')
// (21, 15, 'lutff_0/out')
// (21, 15, 'lutff_2/in_3')
// (21, 16, 'neigh_op_bot_0')
// (22, 14, 'neigh_op_tnl_0')
// (22, 15, 'neigh_op_lft_0')
// (22, 16, 'neigh_op_bnl_0')

wire n1572;
// (20, 14, 'neigh_op_tnr_2')
// (20, 15, 'neigh_op_rgt_2')
// (20, 16, 'neigh_op_bnr_2')
// (21, 14, 'neigh_op_top_2')
// (21, 15, 'lutff_2/out')
// (21, 16, 'local_g1_2')
// (21, 16, 'lutff_7/in_0')
// (21, 16, 'neigh_op_bot_2')
// (22, 14, 'neigh_op_tnl_2')
// (22, 15, 'neigh_op_lft_2')
// (22, 16, 'neigh_op_bnl_2')

wire n1573;
// (20, 14, 'neigh_op_tnr_4')
// (20, 15, 'neigh_op_rgt_4')
// (20, 16, 'neigh_op_bnr_4')
// (21, 14, 'neigh_op_top_4')
// (21, 15, 'lutff_4/out')
// (21, 16, 'neigh_op_bot_4')
// (22, 14, 'neigh_op_tnl_4')
// (22, 15, 'neigh_op_lft_4')
// (22, 16, 'local_g2_4')
// (22, 16, 'lutff_7/in_1')
// (22, 16, 'neigh_op_bnl_4')

reg n1574 = 0;
// (20, 14, 'neigh_op_tnr_5')
// (20, 15, 'neigh_op_rgt_5')
// (20, 16, 'neigh_op_bnr_5')
// (21, 14, 'neigh_op_top_5')
// (21, 15, 'local_g1_5')
// (21, 15, 'lutff_1/in_3')
// (21, 15, 'lutff_5/out')
// (21, 16, 'neigh_op_bot_5')
// (22, 14, 'neigh_op_tnl_5')
// (22, 15, 'neigh_op_lft_5')
// (22, 16, 'neigh_op_bnl_5')

wire n1575;
// (20, 14, 'neigh_op_tnr_6')
// (20, 15, 'neigh_op_rgt_6')
// (20, 16, 'neigh_op_bnr_6')
// (21, 14, 'neigh_op_top_6')
// (21, 15, 'local_g3_6')
// (21, 15, 'lutff_4/in_3')
// (21, 15, 'lutff_6/out')
// (21, 16, 'neigh_op_bot_6')
// (22, 14, 'neigh_op_tnl_6')
// (22, 15, 'neigh_op_lft_6')
// (22, 16, 'neigh_op_bnl_6')

reg n1576 = 0;
// (20, 14, 'neigh_op_tnr_7')
// (20, 15, 'neigh_op_rgt_7')
// (20, 16, 'neigh_op_bnr_7')
// (21, 14, 'neigh_op_top_7')
// (21, 15, 'local_g1_7')
// (21, 15, 'lutff_3/in_3')
// (21, 15, 'lutff_7/out')
// (21, 16, 'neigh_op_bot_7')
// (22, 14, 'neigh_op_tnl_7')
// (22, 15, 'neigh_op_lft_7')
// (22, 16, 'neigh_op_bnl_7')

reg n1577 = 0;
// (20, 14, 'sp4_h_r_10')
// (21, 14, 'local_g0_7')
// (21, 14, 'lutff_6/in_3')
// (21, 14, 'sp4_h_r_23')
// (22, 14, 'sp4_h_r_34')
// (23, 11, 'sp4_r_v_b_40')
// (23, 12, 'neigh_op_tnr_0')
// (23, 12, 'sp4_r_v_b_29')
// (23, 13, 'neigh_op_rgt_0')
// (23, 13, 'sp4_r_v_b_16')
// (23, 14, 'neigh_op_bnr_0')
// (23, 14, 'sp4_h_r_47')
// (23, 14, 'sp4_r_v_b_5')
// (24, 10, 'sp4_v_t_40')
// (24, 11, 'sp4_v_b_40')
// (24, 12, 'neigh_op_top_0')
// (24, 12, 'sp4_v_b_29')
// (24, 13, 'lutff_0/out')
// (24, 13, 'sp4_v_b_16')
// (24, 14, 'neigh_op_bot_0')
// (24, 14, 'sp4_h_l_47')
// (24, 14, 'sp4_v_b_5')
// (25, 12, 'neigh_op_tnl_0')
// (25, 13, 'neigh_op_lft_0')
// (25, 14, 'neigh_op_bnl_0')

wire n1578;
// (20, 15, 'lutff_4/lout')
// (20, 15, 'lutff_5/in_2')

reg n1579 = 0;
// (20, 15, 'neigh_op_tnr_0')
// (20, 16, 'neigh_op_rgt_0')
// (20, 17, 'neigh_op_bnr_0')
// (21, 15, 'neigh_op_top_0')
// (21, 16, 'local_g1_0')
// (21, 16, 'lutff_0/out')
// (21, 16, 'lutff_2/in_3')
// (21, 17, 'neigh_op_bot_0')
// (22, 15, 'neigh_op_tnl_0')
// (22, 16, 'neigh_op_lft_0')
// (22, 17, 'neigh_op_bnl_0')

wire n1580;
// (20, 15, 'neigh_op_tnr_2')
// (20, 16, 'neigh_op_rgt_2')
// (20, 16, 'sp4_r_v_b_36')
// (20, 17, 'neigh_op_bnr_2')
// (20, 17, 'sp4_r_v_b_25')
// (20, 18, 'sp4_r_v_b_12')
// (20, 19, 'sp4_r_v_b_1')
// (21, 15, 'neigh_op_top_2')
// (21, 15, 'sp4_v_t_36')
// (21, 16, 'lutff_2/out')
// (21, 16, 'sp4_v_b_36')
// (21, 17, 'neigh_op_bot_2')
// (21, 17, 'sp4_v_b_25')
// (21, 18, 'sp4_v_b_12')
// (21, 19, 'local_g1_1')
// (21, 19, 'lutff_3/in_1')
// (21, 19, 'sp4_v_b_1')
// (22, 15, 'neigh_op_tnl_2')
// (22, 16, 'neigh_op_lft_2')
// (22, 17, 'neigh_op_bnl_2')

wire n1581;
// (20, 15, 'neigh_op_tnr_4')
// (20, 16, 'neigh_op_rgt_4')
// (20, 17, 'neigh_op_bnr_4')
// (21, 15, 'neigh_op_top_4')
// (21, 16, 'local_g0_4')
// (21, 16, 'lutff_4/out')
// (21, 16, 'lutff_7/in_3')
// (21, 17, 'neigh_op_bot_4')
// (22, 15, 'neigh_op_tnl_4')
// (22, 16, 'neigh_op_lft_4')
// (22, 17, 'neigh_op_bnl_4')

wire n1582;
// (20, 15, 'neigh_op_tnr_7')
// (20, 16, 'neigh_op_rgt_7')
// (20, 17, 'neigh_op_bnr_7')
// (21, 15, 'neigh_op_top_7')
// (21, 16, 'lutff_7/out')
// (21, 17, 'neigh_op_bot_7')
// (22, 15, 'neigh_op_tnl_7')
// (22, 16, 'neigh_op_lft_7')
// (22, 17, 'local_g3_7')
// (22, 17, 'lutff_0/in_0')
// (22, 17, 'neigh_op_bnl_7')

reg n1583 = 0;
// (20, 15, 'sp4_r_v_b_38')
// (20, 16, 'sp4_r_v_b_27')
// (20, 17, 'sp4_r_v_b_14')
// (20, 18, 'sp4_r_v_b_3')
// (21, 14, 'sp4_h_r_3')
// (21, 14, 'sp4_v_t_38')
// (21, 15, 'sp4_v_b_38')
// (21, 16, 'local_g3_3')
// (21, 16, 'lutff_3/in_3')
// (21, 16, 'sp4_v_b_27')
// (21, 17, 'sp4_v_b_14')
// (21, 18, 'sp4_v_b_3')
// (22, 14, 'sp4_h_r_14')
// (23, 13, 'neigh_op_tnr_3')
// (23, 14, 'neigh_op_rgt_3')
// (23, 14, 'sp4_h_r_27')
// (23, 15, 'neigh_op_bnr_3')
// (24, 13, 'neigh_op_top_3')
// (24, 14, 'lutff_3/out')
// (24, 14, 'sp4_h_r_38')
// (24, 15, 'neigh_op_bot_3')
// (25, 13, 'neigh_op_tnl_3')
// (25, 14, 'neigh_op_lft_3')
// (25, 14, 'sp4_h_l_38')
// (25, 15, 'neigh_op_bnl_3')

wire n1584;
// (20, 16, 'neigh_op_tnr_0')
// (20, 17, 'neigh_op_rgt_0')
// (20, 18, 'neigh_op_bnr_0')
// (21, 16, 'neigh_op_top_0')
// (21, 17, 'lutff_0/out')
// (21, 18, 'neigh_op_bot_0')
// (22, 16, 'neigh_op_tnl_0')
// (22, 17, 'local_g0_0')
// (22, 17, 'lutff_3/in_1')
// (22, 17, 'neigh_op_lft_0')
// (22, 18, 'neigh_op_bnl_0')

reg n1585 = 0;
// (20, 16, 'neigh_op_tnr_1')
// (20, 17, 'neigh_op_rgt_1')
// (20, 18, 'neigh_op_bnr_1')
// (21, 16, 'neigh_op_top_1')
// (21, 17, 'local_g2_1')
// (21, 17, 'lutff_0/in_3')
// (21, 17, 'lutff_1/out')
// (21, 18, 'neigh_op_bot_1')
// (22, 16, 'neigh_op_tnl_1')
// (22, 17, 'neigh_op_lft_1')
// (22, 18, 'neigh_op_bnl_1')

wire n1586;
// (20, 16, 'neigh_op_tnr_2')
// (20, 17, 'neigh_op_rgt_2')
// (20, 18, 'neigh_op_bnr_2')
// (21, 16, 'neigh_op_top_2')
// (21, 17, 'lutff_2/out')
// (21, 18, 'neigh_op_bot_2')
// (22, 16, 'neigh_op_tnl_2')
// (22, 17, 'neigh_op_lft_2')
// (22, 18, 'local_g2_2')
// (22, 18, 'lutff_5/in_3')
// (22, 18, 'neigh_op_bnl_2')

reg n1587 = 0;
// (20, 16, 'neigh_op_tnr_3')
// (20, 17, 'neigh_op_rgt_3')
// (20, 18, 'neigh_op_bnr_3')
// (21, 16, 'neigh_op_top_3')
// (21, 17, 'local_g0_3')
// (21, 17, 'lutff_2/in_3')
// (21, 17, 'lutff_3/out')
// (21, 18, 'neigh_op_bot_3')
// (22, 16, 'neigh_op_tnl_3')
// (22, 17, 'neigh_op_lft_3')
// (22, 18, 'neigh_op_bnl_3')

reg n1588 = 0;
// (20, 16, 'neigh_op_tnr_5')
// (20, 17, 'neigh_op_rgt_5')
// (20, 18, 'neigh_op_bnr_5')
// (21, 16, 'neigh_op_top_5')
// (21, 17, 'local_g2_5')
// (21, 17, 'lutff_4/in_3')
// (21, 17, 'lutff_5/out')
// (21, 18, 'neigh_op_bot_5')
// (22, 16, 'neigh_op_tnl_5')
// (22, 17, 'neigh_op_lft_5')
// (22, 18, 'neigh_op_bnl_5')

reg n1589 = 0;
// (20, 16, 'neigh_op_tnr_7')
// (20, 17, 'neigh_op_rgt_7')
// (20, 18, 'neigh_op_bnr_7')
// (21, 16, 'neigh_op_top_7')
// (21, 17, 'local_g2_7')
// (21, 17, 'lutff_6/in_3')
// (21, 17, 'lutff_7/out')
// (21, 18, 'neigh_op_bot_7')
// (22, 16, 'neigh_op_tnl_7')
// (22, 17, 'neigh_op_lft_7')
// (22, 18, 'neigh_op_bnl_7')

reg n1590 = 0;
// (20, 16, 'sp4_h_r_5')
// (21, 16, 'sp4_h_r_16')
// (22, 16, 'local_g3_5')
// (22, 16, 'lutff_5/in_3')
// (22, 16, 'sp4_h_r_29')
// (23, 13, 'neigh_op_tnr_4')
// (23, 13, 'sp4_r_v_b_37')
// (23, 14, 'neigh_op_rgt_4')
// (23, 14, 'sp4_r_v_b_24')
// (23, 15, 'neigh_op_bnr_4')
// (23, 15, 'sp4_r_v_b_13')
// (23, 16, 'sp4_h_r_40')
// (23, 16, 'sp4_r_v_b_0')
// (24, 12, 'sp4_v_t_37')
// (24, 13, 'neigh_op_top_4')
// (24, 13, 'sp4_v_b_37')
// (24, 14, 'lutff_4/out')
// (24, 14, 'sp4_v_b_24')
// (24, 15, 'neigh_op_bot_4')
// (24, 15, 'sp4_v_b_13')
// (24, 16, 'sp4_h_l_40')
// (24, 16, 'sp4_v_b_0')
// (25, 13, 'neigh_op_tnl_4')
// (25, 14, 'neigh_op_lft_4')
// (25, 15, 'neigh_op_bnl_4')

reg n1591 = 0;
// (20, 17, 'local_g1_0')
// (20, 17, 'lutff_0/in_1')
// (20, 17, 'sp12_h_r_0')
// (21, 17, 'sp12_h_r_3')
// (22, 17, 'sp12_h_r_4')
// (23, 16, 'neigh_op_tnr_0')
// (23, 17, 'neigh_op_rgt_0')
// (23, 17, 'sp12_h_r_7')
// (23, 18, 'neigh_op_bnr_0')
// (24, 16, 'neigh_op_top_0')
// (24, 17, 'lutff_0/out')
// (24, 17, 'sp12_h_r_8')
// (24, 18, 'neigh_op_bot_0')
// (25, 16, 'neigh_op_tnl_0')
// (25, 17, 'neigh_op_lft_0')
// (25, 17, 'sp12_h_r_11')
// (25, 18, 'neigh_op_bnl_0')
// (26, 17, 'sp12_h_r_12')
// (27, 17, 'sp12_h_r_15')
// (28, 17, 'sp12_h_r_16')
// (29, 17, 'sp12_h_r_19')
// (30, 17, 'sp12_h_r_20')
// (31, 17, 'sp12_h_r_23')
// (32, 17, 'sp12_h_l_23')

wire n1592;
// (20, 17, 'neigh_op_tnr_1')
// (20, 17, 'sp4_r_v_b_47')
// (20, 18, 'neigh_op_rgt_1')
// (20, 18, 'sp4_r_v_b_34')
// (20, 19, 'neigh_op_bnr_1')
// (20, 19, 'sp4_r_v_b_23')
// (20, 20, 'sp4_r_v_b_10')
// (21, 16, 'sp4_v_t_47')
// (21, 17, 'neigh_op_top_1')
// (21, 17, 'sp4_v_b_47')
// (21, 18, 'lutff_1/out')
// (21, 18, 'sp4_v_b_34')
// (21, 19, 'local_g0_7')
// (21, 19, 'lutff_4/in_1')
// (21, 19, 'neigh_op_bot_1')
// (21, 19, 'sp4_v_b_23')
// (21, 20, 'sp4_v_b_10')
// (22, 17, 'neigh_op_tnl_1')
// (22, 18, 'neigh_op_lft_1')
// (22, 19, 'neigh_op_bnl_1')

reg n1593 = 0;
// (20, 17, 'neigh_op_tnr_2')
// (20, 18, 'neigh_op_rgt_2')
// (20, 19, 'neigh_op_bnr_2')
// (21, 17, 'neigh_op_top_2')
// (21, 18, 'local_g2_2')
// (21, 18, 'lutff_0/in_2')
// (21, 18, 'lutff_2/out')
// (21, 19, 'neigh_op_bot_2')
// (22, 17, 'neigh_op_tnl_2')
// (22, 18, 'neigh_op_lft_2')
// (22, 19, 'neigh_op_bnl_2')

wire n1594;
// (20, 17, 'neigh_op_tnr_4')
// (20, 18, 'neigh_op_rgt_4')
// (20, 19, 'neigh_op_bnr_4')
// (21, 17, 'neigh_op_top_4')
// (21, 18, 'lutff_4/out')
// (21, 19, 'neigh_op_bot_4')
// (22, 17, 'local_g2_4')
// (22, 17, 'lutff_5/in_1')
// (22, 17, 'neigh_op_tnl_4')
// (22, 18, 'neigh_op_lft_4')
// (22, 19, 'neigh_op_bnl_4')

reg n1595 = 0;
// (20, 17, 'neigh_op_tnr_5')
// (20, 18, 'neigh_op_rgt_5')
// (20, 19, 'neigh_op_bnr_5')
// (21, 17, 'neigh_op_top_5')
// (21, 18, 'local_g1_5')
// (21, 18, 'lutff_3/in_3')
// (21, 18, 'lutff_5/out')
// (21, 19, 'neigh_op_bot_5')
// (22, 17, 'neigh_op_tnl_5')
// (22, 18, 'neigh_op_lft_5')
// (22, 19, 'neigh_op_bnl_5')

wire n1596;
// (20, 17, 'neigh_op_tnr_7')
// (20, 18, 'neigh_op_rgt_7')
// (20, 19, 'neigh_op_bnr_7')
// (21, 17, 'neigh_op_top_7')
// (21, 18, 'lutff_7/out')
// (21, 19, 'neigh_op_bot_7')
// (22, 17, 'neigh_op_tnl_7')
// (22, 18, 'local_g1_7')
// (22, 18, 'lutff_0/in_0')
// (22, 18, 'neigh_op_lft_7')
// (22, 19, 'neigh_op_bnl_7')

reg n1597 = 0;
// (20, 17, 'sp4_r_v_b_43')
// (20, 18, 'sp4_r_v_b_30')
// (20, 19, 'sp4_r_v_b_19')
// (20, 20, 'sp4_r_v_b_6')
// (21, 16, 'sp4_h_r_0')
// (21, 16, 'sp4_v_t_43')
// (21, 17, 'local_g2_3')
// (21, 17, 'lutff_2/in_1')
// (21, 17, 'sp4_v_b_43')
// (21, 18, 'sp4_v_b_30')
// (21, 19, 'sp4_v_b_19')
// (21, 20, 'sp4_v_b_6')
// (22, 15, 'neigh_op_tnr_4')
// (22, 16, 'neigh_op_rgt_4')
// (22, 16, 'sp4_h_r_13')
// (22, 17, 'neigh_op_bnr_4')
// (23, 15, 'neigh_op_top_4')
// (23, 16, 'lutff_4/out')
// (23, 16, 'sp4_h_r_24')
// (23, 17, 'neigh_op_bot_4')
// (24, 15, 'neigh_op_tnl_4')
// (24, 16, 'neigh_op_lft_4')
// (24, 16, 'sp4_h_r_37')
// (24, 17, 'neigh_op_bnl_4')
// (25, 16, 'sp4_h_l_37')

reg n1598 = 0;
// (20, 17, 'sp4_r_v_b_45')
// (20, 18, 'sp4_r_v_b_32')
// (20, 19, 'sp4_r_v_b_21')
// (20, 20, 'sp4_r_v_b_8')
// (21, 16, 'sp4_h_r_2')
// (21, 16, 'sp4_v_t_45')
// (21, 17, 'local_g3_5')
// (21, 17, 'lutff_4/in_0')
// (21, 17, 'sp4_v_b_45')
// (21, 18, 'sp4_v_b_32')
// (21, 19, 'sp4_v_b_21')
// (21, 20, 'sp4_v_b_8')
// (22, 15, 'neigh_op_tnr_5')
// (22, 16, 'neigh_op_rgt_5')
// (22, 16, 'sp4_h_r_15')
// (22, 17, 'neigh_op_bnr_5')
// (23, 15, 'neigh_op_top_5')
// (23, 16, 'lutff_5/out')
// (23, 16, 'sp4_h_r_26')
// (23, 17, 'neigh_op_bot_5')
// (24, 15, 'neigh_op_tnl_5')
// (24, 16, 'neigh_op_lft_5')
// (24, 16, 'sp4_h_r_39')
// (24, 17, 'neigh_op_bnl_5')
// (25, 16, 'sp4_h_l_39')

reg n1599 = 0;
// (20, 18, 'local_g3_0')
// (20, 18, 'lutff_0/in_1')
// (20, 18, 'sp4_r_v_b_40')
// (20, 19, 'neigh_op_tnr_0')
// (20, 19, 'sp4_r_v_b_29')
// (20, 20, 'neigh_op_rgt_0')
// (20, 20, 'sp4_r_v_b_16')
// (20, 21, 'neigh_op_bnr_0')
// (20, 21, 'sp4_r_v_b_5')
// (21, 17, 'sp4_v_t_40')
// (21, 18, 'sp4_v_b_40')
// (21, 19, 'neigh_op_top_0')
// (21, 19, 'sp4_v_b_29')
// (21, 20, 'lutff_0/out')
// (21, 20, 'sp4_v_b_16')
// (21, 21, 'neigh_op_bot_0')
// (21, 21, 'sp4_v_b_5')
// (22, 19, 'neigh_op_tnl_0')
// (22, 20, 'neigh_op_lft_0')
// (22, 21, 'neigh_op_bnl_0')

reg n1600 = 0;
// (20, 18, 'local_g3_4')
// (20, 18, 'lutff_5/in_0')
// (20, 18, 'sp4_r_v_b_44')
// (20, 19, 'neigh_op_tnr_2')
// (20, 19, 'sp4_r_v_b_33')
// (20, 20, 'neigh_op_rgt_2')
// (20, 20, 'sp4_r_v_b_20')
// (20, 21, 'neigh_op_bnr_2')
// (20, 21, 'sp4_r_v_b_9')
// (21, 17, 'sp4_v_t_44')
// (21, 18, 'sp4_v_b_44')
// (21, 19, 'neigh_op_top_2')
// (21, 19, 'sp4_v_b_33')
// (21, 20, 'lutff_2/out')
// (21, 20, 'sp4_v_b_20')
// (21, 21, 'neigh_op_bot_2')
// (21, 21, 'sp4_v_b_9')
// (22, 19, 'neigh_op_tnl_2')
// (22, 20, 'neigh_op_lft_2')
// (22, 21, 'neigh_op_bnl_2')

wire n1601;
// (20, 18, 'neigh_op_tnr_2')
// (20, 19, 'neigh_op_rgt_2')
// (20, 20, 'neigh_op_bnr_2')
// (21, 18, 'neigh_op_top_2')
// (21, 19, 'local_g0_2')
// (21, 19, 'lutff_2/out')
// (21, 19, 'lutff_5/in_3')
// (21, 20, 'neigh_op_bot_2')
// (22, 18, 'neigh_op_tnl_2')
// (22, 19, 'neigh_op_lft_2')
// (22, 20, 'neigh_op_bnl_2')

reg n1602 = 0;
// (20, 18, 'sp4_h_r_1')
// (21, 18, 'local_g0_4')
// (21, 18, 'lutff_6/in_2')
// (21, 18, 'sp4_h_r_12')
// (22, 18, 'sp4_h_r_25')
// (23, 14, 'neigh_op_tnr_2')
// (23, 15, 'neigh_op_rgt_2')
// (23, 15, 'sp4_r_v_b_36')
// (23, 16, 'neigh_op_bnr_2')
// (23, 16, 'sp4_r_v_b_25')
// (23, 17, 'sp4_r_v_b_12')
// (23, 18, 'sp4_h_r_36')
// (23, 18, 'sp4_r_v_b_1')
// (24, 14, 'neigh_op_top_2')
// (24, 14, 'sp4_v_t_36')
// (24, 15, 'lutff_2/out')
// (24, 15, 'sp4_v_b_36')
// (24, 16, 'neigh_op_bot_2')
// (24, 16, 'sp4_v_b_25')
// (24, 17, 'sp4_v_b_12')
// (24, 18, 'sp4_h_l_36')
// (24, 18, 'sp4_v_b_1')
// (25, 14, 'neigh_op_tnl_2')
// (25, 15, 'neigh_op_lft_2')
// (25, 16, 'neigh_op_bnl_2')

reg n1603 = 0;
// (20, 19, 'neigh_op_tnr_1')
// (20, 19, 'sp4_r_v_b_47')
// (20, 20, 'neigh_op_rgt_1')
// (20, 20, 'sp4_r_v_b_34')
// (20, 21, 'neigh_op_bnr_1')
// (20, 21, 'sp4_r_v_b_23')
// (20, 22, 'sp4_r_v_b_10')
// (21, 18, 'sp4_v_t_47')
// (21, 19, 'neigh_op_top_1')
// (21, 19, 'sp4_v_b_47')
// (21, 20, 'lutff_1/out')
// (21, 20, 'sp4_v_b_34')
// (21, 21, 'neigh_op_bot_1')
// (21, 21, 'sp4_v_b_23')
// (21, 22, 'local_g1_2')
// (21, 22, 'lutff_2/in_1')
// (21, 22, 'sp4_v_b_10')
// (22, 19, 'neigh_op_tnl_1')
// (22, 20, 'neigh_op_lft_1')
// (22, 21, 'neigh_op_bnl_1')

reg n1604 = 0;
// (20, 19, 'neigh_op_tnr_3')
// (20, 20, 'neigh_op_rgt_3')
// (20, 20, 'sp4_r_v_b_38')
// (20, 21, 'neigh_op_bnr_3')
// (20, 21, 'sp4_r_v_b_27')
// (20, 22, 'sp4_r_v_b_14')
// (20, 23, 'sp4_r_v_b_3')
// (21, 19, 'neigh_op_top_3')
// (21, 19, 'sp4_v_t_38')
// (21, 20, 'lutff_3/out')
// (21, 20, 'sp4_v_b_38')
// (21, 21, 'neigh_op_bot_3')
// (21, 21, 'sp4_v_b_27')
// (21, 22, 'local_g0_6')
// (21, 22, 'lutff_5/in_3')
// (21, 22, 'sp4_v_b_14')
// (21, 23, 'sp4_v_b_3')
// (22, 19, 'neigh_op_tnl_3')
// (22, 20, 'neigh_op_lft_3')
// (22, 21, 'neigh_op_bnl_3')

reg n1605 = 0;
// (20, 19, 'neigh_op_tnr_4')
// (20, 20, 'neigh_op_rgt_4')
// (20, 21, 'neigh_op_bnr_4')
// (21, 19, 'neigh_op_top_4')
// (21, 19, 'sp4_r_v_b_36')
// (21, 20, 'lutff_4/out')
// (21, 20, 'sp4_r_v_b_25')
// (21, 21, 'neigh_op_bot_4')
// (21, 21, 'sp4_r_v_b_12')
// (21, 22, 'local_g1_1')
// (21, 22, 'lutff_1/in_1')
// (21, 22, 'sp4_r_v_b_1')
// (22, 18, 'sp4_v_t_36')
// (22, 19, 'neigh_op_tnl_4')
// (22, 19, 'sp4_v_b_36')
// (22, 20, 'neigh_op_lft_4')
// (22, 20, 'sp4_v_b_25')
// (22, 21, 'neigh_op_bnl_4')
// (22, 21, 'sp4_v_b_12')
// (22, 22, 'sp4_v_b_1')

reg n1606 = 0;
// (20, 19, 'neigh_op_tnr_5')
// (20, 20, 'neigh_op_rgt_5')
// (20, 21, 'neigh_op_bnr_5')
// (21, 19, 'neigh_op_top_5')
// (21, 20, 'lutff_5/out')
// (21, 21, 'neigh_op_bot_5')
// (22, 19, 'local_g3_5')
// (22, 19, 'lutff_2/in_0')
// (22, 19, 'neigh_op_tnl_5')
// (22, 20, 'neigh_op_lft_5')
// (22, 21, 'neigh_op_bnl_5')

reg n1607 = 0;
// (20, 19, 'neigh_op_tnr_6')
// (20, 20, 'neigh_op_rgt_6')
// (20, 21, 'neigh_op_bnr_6')
// (21, 19, 'neigh_op_top_6')
// (21, 20, 'lutff_6/out')
// (21, 21, 'neigh_op_bot_6')
// (22, 19, 'local_g3_6')
// (22, 19, 'lutff_4/in_1')
// (22, 19, 'neigh_op_tnl_6')
// (22, 20, 'neigh_op_lft_6')
// (22, 21, 'neigh_op_bnl_6')

reg n1608 = 0;
// (20, 19, 'sp4_h_r_1')
// (21, 19, 'local_g1_4')
// (21, 19, 'lutff_6/in_1')
// (21, 19, 'sp4_h_r_12')
// (22, 11, 'neigh_op_tnr_2')
// (22, 12, 'neigh_op_rgt_2')
// (22, 13, 'neigh_op_bnr_2')
// (22, 19, 'sp4_h_r_25')
// (23, 11, 'neigh_op_top_2')
// (23, 12, 'lutff_2/out')
// (23, 12, 'sp4_r_v_b_37')
// (23, 13, 'neigh_op_bot_2')
// (23, 13, 'sp4_r_v_b_24')
// (23, 14, 'sp4_r_v_b_13')
// (23, 15, 'sp4_r_v_b_0')
// (23, 16, 'sp4_r_v_b_45')
// (23, 17, 'sp4_r_v_b_32')
// (23, 18, 'sp4_r_v_b_21')
// (23, 19, 'sp4_h_r_36')
// (23, 19, 'sp4_r_v_b_8')
// (24, 11, 'neigh_op_tnl_2')
// (24, 11, 'sp4_v_t_37')
// (24, 12, 'neigh_op_lft_2')
// (24, 12, 'sp4_v_b_37')
// (24, 13, 'neigh_op_bnl_2')
// (24, 13, 'sp4_v_b_24')
// (24, 14, 'sp4_v_b_13')
// (24, 15, 'sp4_v_b_0')
// (24, 15, 'sp4_v_t_45')
// (24, 16, 'sp4_v_b_45')
// (24, 17, 'sp4_v_b_32')
// (24, 18, 'sp4_v_b_21')
// (24, 19, 'sp4_h_l_36')
// (24, 19, 'sp4_v_b_8')

wire n1609;
// (20, 19, 'sp4_r_v_b_39')
// (20, 20, 'sp4_r_v_b_26')
// (20, 21, 'neigh_op_tnr_1')
// (20, 21, 'sp4_r_v_b_15')
// (20, 22, 'neigh_op_rgt_1')
// (20, 22, 'sp4_r_v_b_2')
// (20, 23, 'neigh_op_bnr_1')
// (21, 18, 'sp4_h_r_7')
// (21, 18, 'sp4_v_t_39')
// (21, 19, 'sp4_v_b_39')
// (21, 20, 'sp4_v_b_26')
// (21, 21, 'neigh_op_top_1')
// (21, 21, 'sp4_v_b_15')
// (21, 22, 'lutff_1/out')
// (21, 22, 'sp4_v_b_2')
// (21, 23, 'neigh_op_bot_1')
// (22, 18, 'local_g0_2')
// (22, 18, 'lutff_5/in_1')
// (22, 18, 'sp4_h_r_18')
// (22, 21, 'neigh_op_tnl_1')
// (22, 22, 'neigh_op_lft_1')
// (22, 23, 'neigh_op_bnl_1')
// (23, 18, 'sp4_h_r_31')
// (24, 18, 'sp4_h_r_42')
// (25, 18, 'sp4_h_l_42')

wire n1610;
// (20, 19, 'sp4_r_v_b_43')
// (20, 20, 'sp4_r_v_b_30')
// (20, 21, 'neigh_op_tnr_3')
// (20, 21, 'sp4_r_v_b_19')
// (20, 22, 'neigh_op_rgt_3')
// (20, 22, 'sp4_r_v_b_6')
// (20, 23, 'neigh_op_bnr_3')
// (21, 18, 'sp4_v_t_43')
// (21, 19, 'local_g2_3')
// (21, 19, 'lutff_0/in_3')
// (21, 19, 'sp4_v_b_43')
// (21, 20, 'sp4_v_b_30')
// (21, 21, 'neigh_op_top_3')
// (21, 21, 'sp4_v_b_19')
// (21, 22, 'lutff_3/out')
// (21, 22, 'sp4_v_b_6')
// (21, 23, 'neigh_op_bot_3')
// (22, 21, 'neigh_op_tnl_3')
// (22, 22, 'neigh_op_lft_3')
// (22, 23, 'neigh_op_bnl_3')

wire n1611;
// (20, 20, 'neigh_op_tnr_4')
// (20, 21, 'neigh_op_rgt_4')
// (20, 22, 'neigh_op_bnr_4')
// (21, 20, 'neigh_op_top_4')
// (21, 21, 'local_g1_4')
// (21, 21, 'lutff_2/in_3')
// (21, 21, 'lutff_4/out')
// (21, 22, 'neigh_op_bot_4')
// (22, 20, 'neigh_op_tnl_4')
// (22, 21, 'neigh_op_lft_4')
// (22, 22, 'neigh_op_bnl_4')

wire n1612;
// (20, 20, 'neigh_op_tnr_5')
// (20, 21, 'neigh_op_rgt_5')
// (20, 22, 'neigh_op_bnr_5')
// (21, 20, 'neigh_op_top_5')
// (21, 21, 'local_g2_5')
// (21, 21, 'lutff_2/in_1')
// (21, 21, 'lutff_5/out')
// (21, 22, 'neigh_op_bot_5')
// (22, 20, 'neigh_op_tnl_5')
// (22, 21, 'neigh_op_lft_5')
// (22, 22, 'neigh_op_bnl_5')

reg n1613 = 0;
// (20, 20, 'neigh_op_tnr_6')
// (20, 21, 'neigh_op_rgt_6')
// (20, 22, 'neigh_op_bnr_6')
// (21, 20, 'neigh_op_top_6')
// (21, 21, 'local_g3_6')
// (21, 21, 'lutff_0/in_3')
// (21, 21, 'lutff_6/out')
// (21, 22, 'neigh_op_bot_6')
// (22, 20, 'neigh_op_tnl_6')
// (22, 21, 'neigh_op_lft_6')
// (22, 22, 'neigh_op_bnl_6')

wire n1614;
// (20, 20, 'neigh_op_tnr_7')
// (20, 21, 'neigh_op_rgt_7')
// (20, 22, 'neigh_op_bnr_7')
// (21, 20, 'neigh_op_top_7')
// (21, 21, 'lutff_7/out')
// (21, 22, 'neigh_op_bot_7')
// (22, 20, 'local_g2_7')
// (22, 20, 'lutff_0/in_3')
// (22, 20, 'neigh_op_tnl_7')
// (22, 21, 'neigh_op_lft_7')
// (22, 22, 'neigh_op_bnl_7')

reg n1615 = 0;
// (20, 20, 'sp4_r_v_b_36')
// (20, 21, 'sp4_r_v_b_25')
// (20, 22, 'sp4_r_v_b_12')
// (20, 23, 'sp4_r_v_b_1')
// (21, 18, 'neigh_op_tnr_1')
// (21, 19, 'neigh_op_rgt_1')
// (21, 19, 'sp4_h_r_7')
// (21, 19, 'sp4_v_t_36')
// (21, 20, 'neigh_op_bnr_1')
// (21, 20, 'sp4_v_b_36')
// (21, 21, 'sp4_v_b_25')
// (21, 22, 'local_g0_4')
// (21, 22, 'lutff_1/in_3')
// (21, 22, 'sp4_v_b_12')
// (21, 23, 'sp4_v_b_1')
// (22, 18, 'neigh_op_top_1')
// (22, 19, 'lutff_1/out')
// (22, 19, 'sp4_h_r_18')
// (22, 20, 'neigh_op_bot_1')
// (23, 18, 'neigh_op_tnl_1')
// (23, 19, 'neigh_op_lft_1')
// (23, 19, 'sp4_h_r_31')
// (23, 20, 'neigh_op_bnl_1')
// (24, 19, 'sp4_h_r_42')
// (25, 19, 'sp4_h_l_42')

wire n1616;
// (20, 21, 'neigh_op_tnr_0')
// (20, 22, 'neigh_op_rgt_0')
// (20, 23, 'neigh_op_bnr_0')
// (21, 21, 'local_g0_0')
// (21, 21, 'lutff_7/in_1')
// (21, 21, 'neigh_op_top_0')
// (21, 22, 'lutff_0/out')
// (21, 23, 'neigh_op_bot_0')
// (22, 21, 'neigh_op_tnl_0')
// (22, 22, 'neigh_op_lft_0')
// (22, 23, 'neigh_op_bnl_0')

wire n1617;
// (20, 21, 'neigh_op_tnr_5')
// (20, 22, 'neigh_op_rgt_5')
// (20, 23, 'neigh_op_bnr_5')
// (21, 15, 'sp4_r_v_b_42')
// (21, 16, 'sp4_r_v_b_31')
// (21, 17, 'sp4_r_v_b_18')
// (21, 18, 'sp4_r_v_b_7')
// (21, 19, 'sp4_r_v_b_46')
// (21, 20, 'sp4_r_v_b_35')
// (21, 21, 'neigh_op_top_5')
// (21, 21, 'sp4_r_v_b_22')
// (21, 22, 'lutff_5/out')
// (21, 22, 'sp4_r_v_b_11')
// (21, 23, 'neigh_op_bot_5')
// (22, 14, 'sp4_v_t_42')
// (22, 15, 'sp4_v_b_42')
// (22, 16, 'sp4_v_b_31')
// (22, 17, 'local_g0_2')
// (22, 17, 'lutff_3/in_3')
// (22, 17, 'sp4_v_b_18')
// (22, 18, 'sp4_v_b_7')
// (22, 18, 'sp4_v_t_46')
// (22, 19, 'sp4_v_b_46')
// (22, 20, 'sp4_v_b_35')
// (22, 21, 'neigh_op_tnl_5')
// (22, 21, 'sp4_v_b_22')
// (22, 22, 'neigh_op_lft_5')
// (22, 22, 'sp4_v_b_11')
// (22, 23, 'neigh_op_bnl_5')

wire n1618;
// (20, 22, 'lutff_1/lout')
// (20, 22, 'lutff_2/in_2')

wire n1619;
// (20, 22, 'lutff_3/lout')
// (20, 22, 'lutff_4/in_2')

reg n1620 = 0;
// (20, 23, 'neigh_op_tnr_0')
// (20, 24, 'local_g2_0')
// (20, 24, 'lutff_7/in_1')
// (20, 24, 'neigh_op_rgt_0')
// (20, 25, 'neigh_op_bnr_0')
// (21, 23, 'neigh_op_top_0')
// (21, 24, 'lutff_0/out')
// (21, 25, 'neigh_op_bot_0')
// (22, 23, 'neigh_op_tnl_0')
// (22, 24, 'neigh_op_lft_0')
// (22, 25, 'neigh_op_bnl_0')

reg n1621 = 0;
// (20, 23, 'neigh_op_tnr_1')
// (20, 24, 'local_g0_7')
// (20, 24, 'lutff_7/in_2')
// (20, 24, 'neigh_op_rgt_1')
// (20, 24, 'sp4_h_r_7')
// (20, 25, 'neigh_op_bnr_1')
// (21, 23, 'neigh_op_top_1')
// (21, 24, 'lutff_1/out')
// (21, 24, 'sp4_h_r_18')
// (21, 25, 'neigh_op_bot_1')
// (22, 23, 'neigh_op_tnl_1')
// (22, 24, 'neigh_op_lft_1')
// (22, 24, 'sp4_h_r_31')
// (22, 25, 'neigh_op_bnl_1')
// (23, 24, 'sp4_h_r_42')
// (24, 24, 'sp4_h_l_42')

reg n1622 = 0;
// (21, 9, 'neigh_op_tnr_1')
// (21, 10, 'local_g3_1')
// (21, 10, 'lutff_3/in_3')
// (21, 10, 'neigh_op_rgt_1')
// (21, 11, 'neigh_op_bnr_1')
// (22, 9, 'neigh_op_top_1')
// (22, 10, 'local_g3_1')
// (22, 10, 'lutff_1/in_1')
// (22, 10, 'lutff_1/out')
// (22, 11, 'neigh_op_bot_1')
// (23, 9, 'neigh_op_tnl_1')
// (23, 10, 'neigh_op_lft_1')
// (23, 11, 'neigh_op_bnl_1')

reg n1623 = 0;
// (21, 9, 'neigh_op_tnr_2')
// (21, 10, 'local_g2_2')
// (21, 10, 'lutff_1/in_1')
// (21, 10, 'lutff_5/in_1')
// (21, 10, 'lutff_7/in_1')
// (21, 10, 'neigh_op_rgt_2')
// (21, 11, 'neigh_op_bnr_2')
// (22, 9, 'neigh_op_top_2')
// (22, 10, 'local_g1_2')
// (22, 10, 'lutff_2/in_1')
// (22, 10, 'lutff_2/out')
// (22, 11, 'neigh_op_bot_2')
// (23, 9, 'neigh_op_tnl_2')
// (23, 10, 'neigh_op_lft_2')
// (23, 11, 'neigh_op_bnl_2')

reg n1624 = 0;
// (21, 9, 'neigh_op_tnr_3')
// (21, 10, 'local_g1_3')
// (21, 10, 'lutff_0/in_0')
// (21, 10, 'lutff_4/in_0')
// (21, 10, 'neigh_op_rgt_3')
// (21, 10, 'sp4_h_r_11')
// (21, 11, 'neigh_op_bnr_3')
// (22, 9, 'neigh_op_top_3')
// (22, 10, 'local_g1_3')
// (22, 10, 'lutff_3/in_1')
// (22, 10, 'lutff_3/out')
// (22, 10, 'sp4_h_r_22')
// (22, 11, 'neigh_op_bot_3')
// (23, 9, 'neigh_op_tnl_3')
// (23, 10, 'neigh_op_lft_3')
// (23, 10, 'sp4_h_r_35')
// (23, 11, 'neigh_op_bnl_3')
// (24, 10, 'sp4_h_r_46')
// (25, 10, 'sp4_h_l_46')

wire n1625;
// (21, 9, 'neigh_op_tnr_5')
// (21, 10, 'local_g2_5')
// (21, 10, 'lutff_6/in_3')
// (21, 10, 'neigh_op_rgt_5')
// (21, 11, 'neigh_op_bnr_5')
// (22, 9, 'neigh_op_top_5')
// (22, 10, 'lutff_5/out')
// (22, 11, 'neigh_op_bot_5')
// (23, 9, 'neigh_op_tnl_5')
// (23, 10, 'neigh_op_lft_5')
// (23, 11, 'neigh_op_bnl_5')

reg n1626 = 0;
// (21, 9, 'neigh_op_tnr_6')
// (21, 10, 'local_g3_6')
// (21, 10, 'lutff_3/in_0')
// (21, 10, 'neigh_op_rgt_6')
// (21, 11, 'neigh_op_bnr_6')
// (22, 9, 'neigh_op_top_6')
// (22, 10, 'local_g1_6')
// (22, 10, 'lutff_6/in_1')
// (22, 10, 'lutff_6/out')
// (22, 11, 'neigh_op_bot_6')
// (23, 9, 'neigh_op_tnl_6')
// (23, 10, 'neigh_op_lft_6')
// (23, 11, 'neigh_op_bnl_6')

reg n1627 = 0;
// (21, 10, 'local_g3_0')
// (21, 10, 'lutff_3/in_2')
// (21, 10, 'neigh_op_tnr_0')
// (21, 11, 'neigh_op_rgt_0')
// (21, 12, 'neigh_op_bnr_0')
// (22, 10, 'neigh_op_top_0')
// (22, 11, 'local_g1_0')
// (22, 11, 'lutff_0/in_1')
// (22, 11, 'lutff_0/out')
// (22, 12, 'neigh_op_bot_0')
// (23, 10, 'neigh_op_tnl_0')
// (23, 11, 'neigh_op_lft_0')
// (23, 12, 'neigh_op_bnl_0')

wire n1628;
// (21, 10, 'lutff_0/lout')
// (21, 10, 'lutff_1/in_2')

wire n1629;
// (21, 10, 'lutff_4/lout')
// (21, 10, 'lutff_5/in_2')

wire n1630;
// (21, 10, 'lutff_5/lout')
// (21, 10, 'lutff_6/in_2')

wire n1631;
// (21, 10, 'sp4_r_v_b_38')
// (21, 11, 'local_g1_3')
// (21, 11, 'lutff_global/cen')
// (21, 11, 'sp4_r_v_b_27')
// (21, 12, 'sp4_r_v_b_14')
// (21, 13, 'sp4_r_v_b_3')
// (21, 14, 'neigh_op_tnr_4')
// (21, 14, 'sp4_r_v_b_37')
// (21, 15, 'neigh_op_rgt_4')
// (21, 15, 'sp4_r_v_b_24')
// (21, 16, 'neigh_op_bnr_4')
// (21, 16, 'sp4_r_v_b_13')
// (21, 17, 'sp4_r_v_b_0')
// (22, 9, 'sp4_v_t_38')
// (22, 10, 'sp4_v_b_38')
// (22, 11, 'sp4_v_b_27')
// (22, 12, 'sp4_v_b_14')
// (22, 13, 'sp4_v_b_3')
// (22, 13, 'sp4_v_t_37')
// (22, 14, 'neigh_op_top_4')
// (22, 14, 'sp4_v_b_37')
// (22, 15, 'lutff_4/out')
// (22, 15, 'sp4_v_b_24')
// (22, 16, 'neigh_op_bot_4')
// (22, 16, 'sp4_v_b_13')
// (22, 17, 'sp4_v_b_0')
// (23, 14, 'neigh_op_tnl_4')
// (23, 15, 'neigh_op_lft_4')
// (23, 16, 'neigh_op_bnl_4')

reg n1632 = 0;
// (21, 11, 'neigh_op_tnr_0')
// (21, 11, 'sp4_r_v_b_45')
// (21, 12, 'neigh_op_rgt_0')
// (21, 12, 'sp4_r_v_b_32')
// (21, 13, 'neigh_op_bnr_0')
// (21, 13, 'sp4_r_v_b_21')
// (21, 14, 'local_g2_0')
// (21, 14, 'lutff_0/in_0')
// (21, 14, 'sp4_r_v_b_8')
// (22, 10, 'sp4_v_t_45')
// (22, 11, 'neigh_op_top_0')
// (22, 11, 'sp4_v_b_45')
// (22, 12, 'lutff_0/out')
// (22, 12, 'sp4_v_b_32')
// (22, 13, 'neigh_op_bot_0')
// (22, 13, 'sp4_v_b_21')
// (22, 14, 'sp4_v_b_8')
// (23, 11, 'neigh_op_tnl_0')
// (23, 12, 'neigh_op_lft_0')
// (23, 13, 'neigh_op_bnl_0')

reg n1633 = 0;
// (21, 11, 'neigh_op_tnr_1')
// (21, 11, 'sp4_r_v_b_47')
// (21, 12, 'neigh_op_rgt_1')
// (21, 12, 'sp4_r_v_b_34')
// (21, 13, 'neigh_op_bnr_1')
// (21, 13, 'sp4_r_v_b_23')
// (21, 14, 'local_g2_2')
// (21, 14, 'lutff_3/in_1')
// (21, 14, 'sp4_r_v_b_10')
// (22, 10, 'sp4_v_t_47')
// (22, 11, 'neigh_op_top_1')
// (22, 11, 'sp4_v_b_47')
// (22, 12, 'lutff_1/out')
// (22, 12, 'sp4_v_b_34')
// (22, 13, 'neigh_op_bot_1')
// (22, 13, 'sp4_v_b_23')
// (22, 14, 'sp4_v_b_10')
// (23, 11, 'neigh_op_tnl_1')
// (23, 12, 'neigh_op_lft_1')
// (23, 13, 'neigh_op_bnl_1')

reg n1634 = 0;
// (21, 11, 'neigh_op_tnr_2')
// (21, 12, 'neigh_op_rgt_2')
// (21, 12, 'sp4_r_v_b_36')
// (21, 13, 'neigh_op_bnr_2')
// (21, 13, 'sp4_r_v_b_25')
// (21, 14, 'local_g2_4')
// (21, 14, 'lutff_6/in_0')
// (21, 14, 'sp4_r_v_b_12')
// (21, 15, 'sp4_r_v_b_1')
// (22, 11, 'neigh_op_top_2')
// (22, 11, 'sp4_v_t_36')
// (22, 12, 'lutff_2/out')
// (22, 12, 'sp4_v_b_36')
// (22, 13, 'neigh_op_bot_2')
// (22, 13, 'sp4_v_b_25')
// (22, 14, 'sp4_v_b_12')
// (22, 15, 'sp4_v_b_1')
// (23, 11, 'neigh_op_tnl_2')
// (23, 12, 'neigh_op_lft_2')
// (23, 13, 'neigh_op_bnl_2')

reg n1635 = 0;
// (21, 11, 'neigh_op_tnr_3')
// (21, 12, 'neigh_op_rgt_3')
// (21, 13, 'neigh_op_bnr_3')
// (22, 11, 'neigh_op_top_3')
// (22, 12, 'lutff_3/out')
// (22, 13, 'local_g0_3')
// (22, 13, 'lutff_0/in_1')
// (22, 13, 'neigh_op_bot_3')
// (23, 11, 'neigh_op_tnl_3')
// (23, 12, 'neigh_op_lft_3')
// (23, 13, 'neigh_op_bnl_3')

reg n1636 = 0;
// (21, 11, 'neigh_op_tnr_4')
// (21, 12, 'neigh_op_rgt_4')
// (21, 13, 'neigh_op_bnr_4')
// (22, 11, 'neigh_op_top_4')
// (22, 12, 'lutff_4/out')
// (22, 13, 'local_g0_4')
// (22, 13, 'lutff_3/in_1')
// (22, 13, 'neigh_op_bot_4')
// (23, 11, 'neigh_op_tnl_4')
// (23, 12, 'neigh_op_lft_4')
// (23, 13, 'neigh_op_bnl_4')

reg n1637 = 0;
// (21, 11, 'neigh_op_tnr_5')
// (21, 12, 'neigh_op_rgt_5')
// (21, 13, 'neigh_op_bnr_5')
// (22, 11, 'neigh_op_top_5')
// (22, 12, 'lutff_5/out')
// (22, 13, 'local_g0_5')
// (22, 13, 'lutff_6/in_1')
// (22, 13, 'neigh_op_bot_5')
// (23, 11, 'neigh_op_tnl_5')
// (23, 12, 'neigh_op_lft_5')
// (23, 13, 'neigh_op_bnl_5')

wire n1638;
// (21, 12, 'neigh_op_tnr_1')
// (21, 13, 'neigh_op_rgt_1')
// (21, 14, 'neigh_op_bnr_1')
// (22, 10, 'sp12_v_t_22')
// (22, 11, 'sp12_v_b_22')
// (22, 12, 'neigh_op_top_1')
// (22, 12, 'sp12_v_b_21')
// (22, 13, 'lutff_1/out')
// (22, 13, 'sp12_v_b_18')
// (22, 14, 'neigh_op_bot_1')
// (22, 14, 'sp12_v_b_17')
// (22, 15, 'sp12_v_b_14')
// (22, 16, 'sp12_v_b_13')
// (22, 17, 'local_g2_2')
// (22, 17, 'lutff_5/in_3')
// (22, 17, 'sp12_v_b_10')
// (22, 18, 'sp12_v_b_9')
// (22, 19, 'sp12_v_b_6')
// (22, 20, 'sp12_v_b_5')
// (22, 21, 'sp12_v_b_2')
// (22, 22, 'sp12_v_b_1')
// (23, 12, 'neigh_op_tnl_1')
// (23, 13, 'neigh_op_lft_1')
// (23, 14, 'neigh_op_bnl_1')

reg n1639 = 0;
// (21, 12, 'neigh_op_tnr_2')
// (21, 13, 'neigh_op_rgt_2')
// (21, 14, 'neigh_op_bnr_2')
// (22, 12, 'neigh_op_top_2')
// (22, 13, 'local_g3_2')
// (22, 13, 'lutff_0/in_3')
// (22, 13, 'lutff_2/out')
// (22, 14, 'neigh_op_bot_2')
// (23, 12, 'neigh_op_tnl_2')
// (23, 13, 'neigh_op_lft_2')
// (23, 14, 'neigh_op_bnl_2')

wire n1640;
// (21, 12, 'neigh_op_tnr_4')
// (21, 13, 'neigh_op_rgt_4')
// (21, 13, 'sp4_r_v_b_40')
// (21, 14, 'neigh_op_bnr_4')
// (21, 14, 'sp4_r_v_b_29')
// (21, 15, 'sp4_r_v_b_16')
// (21, 16, 'sp4_r_v_b_5')
// (21, 17, 'sp4_r_v_b_40')
// (21, 18, 'sp4_r_v_b_29')
// (21, 19, 'sp4_r_v_b_16')
// (21, 20, 'sp4_r_v_b_5')
// (22, 12, 'neigh_op_top_4')
// (22, 12, 'sp4_v_t_40')
// (22, 13, 'lutff_4/out')
// (22, 13, 'sp4_v_b_40')
// (22, 14, 'neigh_op_bot_4')
// (22, 14, 'sp4_v_b_29')
// (22, 15, 'sp4_v_b_16')
// (22, 16, 'sp4_v_b_5')
// (22, 16, 'sp4_v_t_40')
// (22, 17, 'sp4_v_b_40')
// (22, 18, 'local_g2_5')
// (22, 18, 'lutff_0/in_1')
// (22, 18, 'sp4_v_b_29')
// (22, 19, 'sp4_v_b_16')
// (22, 20, 'sp4_v_b_5')
// (23, 12, 'neigh_op_tnl_4')
// (23, 13, 'neigh_op_lft_4')
// (23, 14, 'neigh_op_bnl_4')

reg n1641 = 0;
// (21, 12, 'neigh_op_tnr_5')
// (21, 13, 'neigh_op_rgt_5')
// (21, 14, 'neigh_op_bnr_5')
// (22, 12, 'neigh_op_top_5')
// (22, 13, 'local_g1_5')
// (22, 13, 'lutff_3/in_3')
// (22, 13, 'lutff_5/out')
// (22, 14, 'neigh_op_bot_5')
// (23, 12, 'neigh_op_tnl_5')
// (23, 13, 'neigh_op_lft_5')
// (23, 14, 'neigh_op_bnl_5')

reg n1642 = 0;
// (21, 13, 'local_g3_1')
// (21, 13, 'lutff_7/in_3')
// (21, 13, 'neigh_op_tnr_1')
// (21, 14, 'neigh_op_rgt_1')
// (21, 15, 'neigh_op_bnr_1')
// (22, 13, 'neigh_op_top_1')
// (22, 14, 'lutff_1/out')
// (22, 15, 'neigh_op_bot_1')
// (23, 13, 'neigh_op_tnl_1')
// (23, 14, 'neigh_op_lft_1')
// (23, 15, 'neigh_op_bnl_1')

wire n1643;
// (21, 13, 'lutff_1/lout')
// (21, 13, 'lutff_2/in_2')

wire n1644;
// (21, 13, 'lutff_2/lout')
// (21, 13, 'lutff_3/in_2')

wire n1645;
// (21, 13, 'lutff_5/lout')
// (21, 13, 'lutff_6/in_2')

reg n1646 = 0;
// (21, 13, 'neigh_op_tnr_2')
// (21, 14, 'neigh_op_rgt_2')
// (21, 14, 'sp4_r_v_b_36')
// (21, 15, 'neigh_op_bnr_2')
// (21, 15, 'sp4_r_v_b_25')
// (21, 16, 'local_g2_4')
// (21, 16, 'lutff_1/in_3')
// (21, 16, 'sp4_r_v_b_12')
// (21, 17, 'sp4_r_v_b_1')
// (22, 13, 'neigh_op_top_2')
// (22, 13, 'sp4_v_t_36')
// (22, 14, 'lutff_2/out')
// (22, 14, 'sp4_v_b_36')
// (22, 15, 'neigh_op_bot_2')
// (22, 15, 'sp4_v_b_25')
// (22, 16, 'sp4_v_b_12')
// (22, 17, 'sp4_v_b_1')
// (23, 13, 'neigh_op_tnl_2')
// (23, 14, 'neigh_op_lft_2')
// (23, 15, 'neigh_op_bnl_2')

reg n1647 = 0;
// (21, 13, 'neigh_op_tnr_3')
// (21, 14, 'neigh_op_rgt_3')
// (21, 14, 'sp4_r_v_b_38')
// (21, 15, 'neigh_op_bnr_3')
// (21, 15, 'sp4_r_v_b_27')
// (21, 16, 'sp4_r_v_b_14')
// (21, 17, 'sp4_r_v_b_3')
// (22, 13, 'neigh_op_top_3')
// (22, 13, 'sp4_v_t_38')
// (22, 14, 'lutff_3/out')
// (22, 14, 'sp4_v_b_38')
// (22, 15, 'neigh_op_bot_3')
// (22, 15, 'sp4_v_b_27')
// (22, 16, 'local_g0_6')
// (22, 16, 'lutff_1/in_3')
// (22, 16, 'sp4_v_b_14')
// (22, 17, 'sp4_v_b_3')
// (23, 13, 'neigh_op_tnl_3')
// (23, 14, 'neigh_op_lft_3')
// (23, 15, 'neigh_op_bnl_3')

wire n1648;
// (21, 14, 'lutff_0/lout')
// (21, 14, 'lutff_1/in_2')

wire n1649;
// (21, 14, 'lutff_3/lout')
// (21, 14, 'lutff_4/in_2')

wire n1650;
// (21, 14, 'lutff_6/lout')
// (21, 14, 'lutff_7/in_2')

wire n1651;
// (21, 14, 'neigh_op_tnr_0')
// (21, 15, 'neigh_op_rgt_0')
// (21, 16, 'neigh_op_bnr_0')
// (22, 11, 'sp12_v_t_23')
// (22, 12, 'sp12_v_b_23')
// (22, 13, 'sp12_v_b_20')
// (22, 14, 'local_g3_3')
// (22, 14, 'lutff_global/cen')
// (22, 14, 'neigh_op_top_0')
// (22, 14, 'sp12_v_b_19')
// (22, 15, 'lutff_0/out')
// (22, 15, 'sp12_v_b_16')
// (22, 16, 'neigh_op_bot_0')
// (22, 16, 'sp12_v_b_15')
// (22, 17, 'sp12_v_b_12')
// (22, 18, 'sp12_v_b_11')
// (22, 19, 'sp12_v_b_8')
// (22, 20, 'sp12_v_b_7')
// (22, 21, 'sp12_v_b_4')
// (22, 22, 'sp12_v_b_3')
// (22, 23, 'sp12_v_b_0')
// (23, 14, 'neigh_op_tnl_0')
// (23, 15, 'neigh_op_lft_0')
// (23, 16, 'neigh_op_bnl_0')

wire n1652;
// (21, 14, 'neigh_op_tnr_1')
// (21, 14, 'sp4_r_v_b_47')
// (21, 15, 'neigh_op_rgt_1')
// (21, 15, 'sp4_r_v_b_34')
// (21, 16, 'neigh_op_bnr_1')
// (21, 16, 'sp4_r_v_b_23')
// (21, 17, 'sp4_r_v_b_10')
// (21, 18, 'sp4_r_v_b_47')
// (21, 19, 'sp4_r_v_b_34')
// (21, 20, 'sp4_r_v_b_23')
// (21, 21, 'sp4_r_v_b_10')
// (22, 13, 'sp4_v_t_47')
// (22, 14, 'neigh_op_top_1')
// (22, 14, 'sp4_v_b_47')
// (22, 15, 'lutff_1/out')
// (22, 15, 'sp4_v_b_34')
// (22, 16, 'neigh_op_bot_1')
// (22, 16, 'sp4_v_b_23')
// (22, 17, 'sp4_v_b_10')
// (22, 17, 'sp4_v_t_47')
// (22, 18, 'sp4_v_b_47')
// (22, 19, 'sp4_v_b_34')
// (22, 20, 'sp4_v_b_23')
// (22, 21, 'local_g0_2')
// (22, 21, 'lutff_global/cen')
// (22, 21, 'sp4_v_b_10')
// (23, 14, 'neigh_op_tnl_1')
// (23, 15, 'neigh_op_lft_1')
// (23, 16, 'neigh_op_bnl_1')

wire n1653;
// (21, 14, 'neigh_op_tnr_3')
// (21, 15, 'neigh_op_rgt_3')
// (21, 16, 'neigh_op_bnr_3')
// (22, 14, 'neigh_op_top_3')
// (22, 15, 'lutff_3/out')
// (22, 16, 'neigh_op_bot_3')
// (23, 14, 'neigh_op_tnl_3')
// (23, 15, 'neigh_op_lft_3')
// (23, 16, 'local_g3_3')
// (23, 16, 'lutff_global/cen')
// (23, 16, 'neigh_op_bnl_3')

wire n1654;
// (21, 14, 'neigh_op_tnr_5')
// (21, 15, 'neigh_op_rgt_5')
// (21, 16, 'neigh_op_bnr_5')
// (22, 14, 'neigh_op_top_5')
// (22, 15, 'lutff_5/out')
// (22, 15, 'sp4_r_v_b_43')
// (22, 16, 'neigh_op_bot_5')
// (22, 16, 'sp4_r_v_b_30')
// (22, 17, 'sp4_r_v_b_19')
// (22, 18, 'sp4_r_v_b_6')
// (23, 14, 'neigh_op_tnl_5')
// (23, 14, 'sp4_v_t_43')
// (23, 15, 'local_g3_3')
// (23, 15, 'lutff_global/cen')
// (23, 15, 'neigh_op_lft_5')
// (23, 15, 'sp4_v_b_43')
// (23, 16, 'neigh_op_bnl_5')
// (23, 16, 'sp4_v_b_30')
// (23, 17, 'sp4_v_b_19')
// (23, 18, 'sp4_v_b_6')

wire n1655;
// (21, 14, 'neigh_op_tnr_6')
// (21, 15, 'neigh_op_rgt_6')
// (21, 16, 'neigh_op_bnr_6')
// (22, 14, 'neigh_op_top_6')
// (22, 15, 'lutff_6/out')
// (22, 15, 'sp4_r_v_b_45')
// (22, 16, 'neigh_op_bot_6')
// (22, 16, 'sp4_r_v_b_32')
// (22, 17, 'sp4_r_v_b_21')
// (22, 18, 'sp4_r_v_b_8')
// (22, 19, 'sp4_r_v_b_46')
// (22, 20, 'sp4_r_v_b_35')
// (22, 21, 'sp4_r_v_b_22')
// (22, 22, 'sp4_r_v_b_11')
// (23, 14, 'neigh_op_tnl_6')
// (23, 14, 'sp4_v_t_45')
// (23, 15, 'neigh_op_lft_6')
// (23, 15, 'sp4_v_b_45')
// (23, 16, 'neigh_op_bnl_6')
// (23, 16, 'sp4_v_b_32')
// (23, 17, 'sp4_v_b_21')
// (23, 18, 'sp4_v_b_8')
// (23, 18, 'sp4_v_t_46')
// (23, 19, 'sp4_v_b_46')
// (23, 20, 'local_g3_3')
// (23, 20, 'lutff_global/cen')
// (23, 20, 'sp4_v_b_35')
// (23, 21, 'sp4_v_b_22')
// (23, 22, 'sp4_v_b_11')

wire n1656;
// (21, 14, 'neigh_op_tnr_7')
// (21, 15, 'neigh_op_rgt_7')
// (21, 16, 'neigh_op_bnr_7')
// (22, 14, 'neigh_op_top_7')
// (22, 15, 'lutff_7/out')
// (22, 15, 'sp4_r_v_b_47')
// (22, 16, 'neigh_op_bot_7')
// (22, 16, 'sp4_r_v_b_34')
// (22, 17, 'sp4_r_v_b_23')
// (22, 18, 'sp4_r_v_b_10')
// (22, 19, 'sp4_r_v_b_43')
// (22, 20, 'sp4_r_v_b_30')
// (22, 21, 'sp4_r_v_b_19')
// (22, 22, 'sp4_r_v_b_6')
// (22, 23, 'local_g3_3')
// (22, 23, 'lutff_global/cen')
// (22, 23, 'sp4_r_v_b_43')
// (22, 24, 'sp4_r_v_b_30')
// (22, 25, 'sp4_r_v_b_19')
// (22, 26, 'sp4_r_v_b_6')
// (23, 14, 'neigh_op_tnl_7')
// (23, 14, 'sp4_v_t_47')
// (23, 15, 'neigh_op_lft_7')
// (23, 15, 'sp4_v_b_47')
// (23, 16, 'neigh_op_bnl_7')
// (23, 16, 'sp4_v_b_34')
// (23, 17, 'sp4_v_b_23')
// (23, 18, 'sp4_v_b_10')
// (23, 18, 'sp4_v_t_43')
// (23, 19, 'sp4_v_b_43')
// (23, 20, 'sp4_v_b_30')
// (23, 21, 'sp4_v_b_19')
// (23, 22, 'sp4_v_b_6')
// (23, 22, 'sp4_v_t_43')
// (23, 23, 'sp4_v_b_43')
// (23, 24, 'sp4_v_b_30')
// (23, 25, 'sp4_v_b_19')
// (23, 26, 'sp4_v_b_6')

wire n1657;
// (21, 15, 'lutff_1/lout')
// (21, 15, 'lutff_2/in_2')

wire n1658;
// (21, 15, 'lutff_3/lout')
// (21, 15, 'lutff_4/in_2')

reg n1659 = 0;
// (21, 15, 'neigh_op_tnr_0')
// (21, 16, 'neigh_op_rgt_0')
// (21, 17, 'neigh_op_bnr_0')
// (22, 15, 'neigh_op_top_0')
// (22, 16, 'local_g1_0')
// (22, 16, 'lutff_0/out')
// (22, 16, 'lutff_2/in_3')
// (22, 17, 'neigh_op_bot_0')
// (23, 15, 'neigh_op_tnl_0')
// (23, 16, 'neigh_op_lft_0')
// (23, 17, 'neigh_op_bnl_0')

wire n1660;
// (21, 15, 'neigh_op_tnr_2')
// (21, 16, 'neigh_op_rgt_2')
// (21, 17, 'neigh_op_bnr_2')
// (22, 15, 'neigh_op_top_2')
// (22, 16, 'lutff_2/out')
// (22, 17, 'local_g1_2')
// (22, 17, 'lutff_4/in_1')
// (22, 17, 'neigh_op_bot_2')
// (23, 15, 'neigh_op_tnl_2')
// (23, 16, 'neigh_op_lft_2')
// (23, 17, 'neigh_op_bnl_2')

wire n1661;
// (21, 15, 'neigh_op_tnr_4')
// (21, 16, 'neigh_op_rgt_4')
// (21, 17, 'neigh_op_bnr_4')
// (22, 15, 'neigh_op_top_4')
// (22, 16, 'local_g0_4')
// (22, 16, 'lutff_4/out')
// (22, 16, 'lutff_7/in_3')
// (22, 17, 'neigh_op_bot_4')
// (23, 15, 'neigh_op_tnl_4')
// (23, 16, 'neigh_op_lft_4')
// (23, 17, 'neigh_op_bnl_4')

wire n1662;
// (21, 15, 'neigh_op_tnr_7')
// (21, 16, 'neigh_op_rgt_7')
// (21, 16, 'sp4_r_v_b_46')
// (21, 17, 'neigh_op_bnr_7')
// (21, 17, 'sp4_r_v_b_35')
// (21, 18, 'sp4_r_v_b_22')
// (21, 19, 'sp4_r_v_b_11')
// (22, 15, 'neigh_op_top_7')
// (22, 15, 'sp4_v_t_46')
// (22, 16, 'lutff_7/out')
// (22, 16, 'sp4_v_b_46')
// (22, 17, 'neigh_op_bot_7')
// (22, 17, 'sp4_v_b_35')
// (22, 18, 'local_g0_6')
// (22, 18, 'lutff_1/in_1')
// (22, 18, 'sp4_v_b_22')
// (22, 19, 'sp4_v_b_11')
// (23, 15, 'neigh_op_tnl_7')
// (23, 16, 'neigh_op_lft_7')
// (23, 17, 'neigh_op_bnl_7')

wire n1663;
// (21, 16, 'lutff_1/lout')
// (21, 16, 'lutff_2/in_2')

wire n1664;
// (21, 16, 'lutff_3/lout')
// (21, 16, 'lutff_4/in_2')

wire n1665;
// (21, 16, 'lutff_5/lout')
// (21, 16, 'lutff_6/in_2')

wire n1666;
// (21, 16, 'lutff_6/lout')
// (21, 16, 'lutff_7/in_2')

wire n1667;
// (21, 16, 'neigh_op_tnr_3')
// (21, 17, 'neigh_op_rgt_3')
// (21, 18, 'neigh_op_bnr_3')
// (22, 16, 'neigh_op_top_3')
// (22, 17, 'local_g0_3')
// (22, 17, 'lutff_3/out')
// (22, 17, 'lutff_6/in_3')
// (22, 18, 'neigh_op_bot_3')
// (23, 16, 'neigh_op_tnl_3')
// (23, 17, 'neigh_op_lft_3')
// (23, 18, 'neigh_op_bnl_3')

wire n1668;
// (21, 16, 'neigh_op_tnr_5')
// (21, 17, 'neigh_op_rgt_5')
// (21, 18, 'neigh_op_bnr_5')
// (22, 16, 'neigh_op_top_5')
// (22, 17, 'local_g0_5')
// (22, 17, 'lutff_0/in_1')
// (22, 17, 'lutff_5/out')
// (22, 18, 'neigh_op_bot_5')
// (23, 16, 'neigh_op_tnl_5')
// (23, 17, 'neigh_op_lft_5')
// (23, 18, 'neigh_op_bnl_5')

wire n1669;
// (21, 16, 'neigh_op_tnr_6')
// (21, 17, 'neigh_op_rgt_6')
// (21, 18, 'neigh_op_bnr_6')
// (22, 16, 'neigh_op_top_6')
// (22, 17, 'local_g3_6')
// (22, 17, 'lutff_0/in_3')
// (22, 17, 'lutff_6/out')
// (22, 18, 'neigh_op_bot_6')
// (23, 16, 'neigh_op_tnl_6')
// (23, 17, 'neigh_op_lft_6')
// (23, 18, 'neigh_op_bnl_6')

wire n1670;
// (21, 17, 'neigh_op_tnr_3')
// (21, 18, 'neigh_op_rgt_3')
// (21, 19, 'neigh_op_bnr_3')
// (22, 17, 'neigh_op_top_3')
// (22, 18, 'local_g0_3')
// (22, 18, 'lutff_0/in_3')
// (22, 18, 'lutff_3/out')
// (22, 19, 'neigh_op_bot_3')
// (23, 17, 'neigh_op_tnl_3')
// (23, 18, 'neigh_op_lft_3')
// (23, 19, 'neigh_op_bnl_3')

wire n1671;
// (21, 17, 'neigh_op_tnr_6')
// (21, 18, 'neigh_op_rgt_6')
// (21, 19, 'neigh_op_bnr_6')
// (22, 17, 'neigh_op_top_6')
// (22, 18, 'local_g2_6')
// (22, 18, 'lutff_1/in_3')
// (22, 18, 'lutff_6/out')
// (22, 19, 'neigh_op_bot_6')
// (23, 17, 'neigh_op_tnl_6')
// (23, 18, 'neigh_op_lft_6')
// (23, 19, 'neigh_op_bnl_6')

wire n1672;
// (21, 17, 'sp4_r_v_b_45')
// (21, 18, 'sp4_r_v_b_32')
// (21, 19, 'neigh_op_tnr_4')
// (21, 19, 'sp4_r_v_b_21')
// (21, 20, 'neigh_op_rgt_4')
// (21, 20, 'sp4_r_v_b_8')
// (21, 21, 'neigh_op_bnr_4')
// (22, 16, 'sp4_v_t_45')
// (22, 17, 'local_g3_5')
// (22, 17, 'lutff_6/in_0')
// (22, 17, 'sp4_v_b_45')
// (22, 18, 'sp4_v_b_32')
// (22, 19, 'neigh_op_top_4')
// (22, 19, 'sp4_v_b_21')
// (22, 20, 'lutff_4/out')
// (22, 20, 'sp4_v_b_8')
// (22, 21, 'neigh_op_bot_4')
// (23, 19, 'neigh_op_tnl_4')
// (23, 20, 'neigh_op_lft_4')
// (23, 21, 'neigh_op_bnl_4')

wire n1673;
// (21, 18, 'lutff_0/lout')
// (21, 18, 'lutff_1/in_2')

wire n1674;
// (21, 18, 'lutff_3/lout')
// (21, 18, 'lutff_4/in_2')

wire n1675;
// (21, 18, 'lutff_6/lout')
// (21, 18, 'lutff_7/in_2')

reg n1676 = 0;
// (21, 18, 'neigh_op_tnr_3')
// (21, 19, 'neigh_op_rgt_3')
// (21, 20, 'neigh_op_bnr_3')
// (22, 18, 'neigh_op_top_3')
// (22, 19, 'local_g0_3')
// (22, 19, 'lutff_2/in_3')
// (22, 19, 'lutff_3/out')
// (22, 20, 'neigh_op_bot_3')
// (23, 18, 'neigh_op_tnl_3')
// (23, 19, 'neigh_op_lft_3')
// (23, 20, 'neigh_op_bnl_3')

reg n1677 = 0;
// (21, 18, 'neigh_op_tnr_5')
// (21, 19, 'neigh_op_rgt_5')
// (21, 20, 'neigh_op_bnr_5')
// (22, 18, 'neigh_op_top_5')
// (22, 19, 'local_g2_5')
// (22, 19, 'lutff_4/in_3')
// (22, 19, 'lutff_5/out')
// (22, 20, 'neigh_op_bot_5')
// (23, 18, 'neigh_op_tnl_5')
// (23, 19, 'neigh_op_lft_5')
// (23, 20, 'neigh_op_bnl_5')

wire n1678;
// (21, 18, 'neigh_op_tnr_7')
// (21, 19, 'neigh_op_rgt_7')
// (21, 20, 'neigh_op_bnr_7')
// (22, 18, 'neigh_op_top_7')
// (22, 19, 'lutff_7/out')
// (22, 20, 'local_g0_7')
// (22, 20, 'lutff_4/in_3')
// (22, 20, 'neigh_op_bot_7')
// (23, 18, 'neigh_op_tnl_7')
// (23, 19, 'neigh_op_lft_7')
// (23, 20, 'neigh_op_bnl_7')

wire n1679;
// (21, 19, 'local_g3_0')
// (21, 19, 'lutff_2/in_3')
// (21, 19, 'neigh_op_tnr_0')
// (21, 20, 'neigh_op_rgt_0')
// (21, 21, 'neigh_op_bnr_0')
// (22, 19, 'neigh_op_top_0')
// (22, 20, 'lutff_0/out')
// (22, 21, 'neigh_op_bot_0')
// (23, 19, 'neigh_op_tnl_0')
// (23, 20, 'neigh_op_lft_0')
// (23, 21, 'neigh_op_bnl_0')

wire n1680;
// (21, 19, 'lutff_0/lout')
// (21, 19, 'lutff_1/in_2')

wire n1681;
// (21, 19, 'lutff_1/lout')
// (21, 19, 'lutff_2/in_2')

wire n1682;
// (21, 19, 'lutff_3/lout')
// (21, 19, 'lutff_4/in_2')

wire n1683;
// (21, 19, 'lutff_4/lout')
// (21, 19, 'lutff_5/in_2')

wire n1684;
// (21, 19, 'lutff_5/lout')
// (21, 19, 'lutff_6/in_2')

wire n1685;
// (21, 19, 'neigh_op_tnr_1')
// (21, 20, 'neigh_op_rgt_1')
// (21, 21, 'neigh_op_bnr_1')
// (22, 19, 'neigh_op_top_1')
// (22, 20, 'local_g2_1')
// (22, 20, 'lutff_0/in_1')
// (22, 20, 'lutff_1/out')
// (22, 21, 'neigh_op_bot_1')
// (23, 19, 'neigh_op_tnl_1')
// (23, 20, 'neigh_op_lft_1')
// (23, 21, 'neigh_op_bnl_1')

reg n1686 = 0;
// (21, 19, 'neigh_op_tnr_5')
// (21, 20, 'neigh_op_rgt_5')
// (21, 21, 'neigh_op_bnr_5')
// (22, 19, 'neigh_op_top_5')
// (22, 20, 'local_g1_5')
// (22, 20, 'lutff_1/in_3')
// (22, 20, 'lutff_5/out')
// (22, 21, 'neigh_op_bot_5')
// (23, 19, 'neigh_op_tnl_5')
// (23, 20, 'neigh_op_lft_5')
// (23, 21, 'neigh_op_bnl_5')

wire n1687;
// (21, 19, 'neigh_op_tnr_6')
// (21, 20, 'neigh_op_rgt_6')
// (21, 21, 'neigh_op_bnr_6')
// (22, 19, 'neigh_op_top_6')
// (22, 20, 'local_g2_6')
// (22, 20, 'lutff_3/in_3')
// (22, 20, 'lutff_6/out')
// (22, 21, 'neigh_op_bot_6')
// (23, 19, 'neigh_op_tnl_6')
// (23, 20, 'neigh_op_lft_6')
// (23, 21, 'neigh_op_bnl_6')

wire n1688;
// (21, 19, 'neigh_op_tnr_7')
// (21, 20, 'neigh_op_rgt_7')
// (21, 21, 'neigh_op_bnr_7')
// (22, 19, 'neigh_op_top_7')
// (22, 20, 'local_g1_7')
// (22, 20, 'lutff_0/in_0')
// (22, 20, 'lutff_7/out')
// (22, 21, 'neigh_op_bot_7')
// (23, 19, 'neigh_op_tnl_7')
// (23, 20, 'neigh_op_lft_7')
// (23, 21, 'neigh_op_bnl_7')

reg n1689 = 0;
// (21, 19, 'sp4_r_v_b_40')
// (21, 20, 'neigh_op_tnr_0')
// (21, 20, 'sp4_r_v_b_29')
// (21, 21, 'neigh_op_rgt_0')
// (21, 21, 'sp4_r_v_b_16')
// (21, 22, 'neigh_op_bnr_0')
// (21, 22, 'sp4_r_v_b_5')
// (22, 18, 'sp4_v_t_40')
// (22, 19, 'local_g3_0')
// (22, 19, 'lutff_6/in_1')
// (22, 19, 'sp4_v_b_40')
// (22, 20, 'neigh_op_top_0')
// (22, 20, 'sp4_v_b_29')
// (22, 21, 'lutff_0/out')
// (22, 21, 'sp4_v_b_16')
// (22, 22, 'neigh_op_bot_0')
// (22, 22, 'sp4_v_b_5')
// (23, 20, 'neigh_op_tnl_0')
// (23, 21, 'neigh_op_lft_0')
// (23, 22, 'neigh_op_bnl_0')

reg n1690 = 0;
// (21, 19, 'sp4_r_v_b_42')
// (21, 20, 'sp4_r_v_b_31')
// (21, 21, 'local_g3_2')
// (21, 21, 'lutff_4/in_3')
// (21, 21, 'sp4_r_v_b_18')
// (21, 22, 'sp4_r_v_b_7')
// (22, 17, 'neigh_op_tnr_1')
// (22, 18, 'neigh_op_rgt_1')
// (22, 18, 'sp4_h_r_7')
// (22, 18, 'sp4_v_t_42')
// (22, 19, 'neigh_op_bnr_1')
// (22, 19, 'sp4_v_b_42')
// (22, 20, 'sp4_v_b_31')
// (22, 21, 'sp4_v_b_18')
// (22, 22, 'sp4_v_b_7')
// (23, 17, 'neigh_op_top_1')
// (23, 18, 'lutff_1/out')
// (23, 18, 'sp4_h_r_18')
// (23, 19, 'neigh_op_bot_1')
// (24, 17, 'neigh_op_tnl_1')
// (24, 18, 'neigh_op_lft_1')
// (24, 18, 'sp4_h_r_31')
// (24, 19, 'neigh_op_bnl_1')
// (25, 18, 'sp4_h_r_42')
// (26, 18, 'sp4_h_l_42')

reg n1691 = 0;
// (21, 20, 'neigh_op_tnr_1')
// (21, 21, 'local_g3_1')
// (21, 21, 'lutff_4/in_0')
// (21, 21, 'neigh_op_rgt_1')
// (21, 22, 'neigh_op_bnr_1')
// (22, 20, 'neigh_op_top_1')
// (22, 21, 'lutff_1/out')
// (22, 22, 'neigh_op_bot_1')
// (23, 20, 'neigh_op_tnl_1')
// (23, 21, 'neigh_op_lft_1')
// (23, 22, 'neigh_op_bnl_1')

reg n1692 = 0;
// (21, 20, 'neigh_op_tnr_2')
// (21, 21, 'neigh_op_rgt_2')
// (21, 22, 'neigh_op_bnr_2')
// (22, 20, 'local_g0_2')
// (22, 20, 'lutff_1/in_1')
// (22, 20, 'neigh_op_top_2')
// (22, 21, 'lutff_2/out')
// (22, 22, 'neigh_op_bot_2')
// (23, 20, 'neigh_op_tnl_2')
// (23, 21, 'neigh_op_lft_2')
// (23, 22, 'neigh_op_bnl_2')

reg n1693 = 0;
// (21, 20, 'neigh_op_tnr_3')
// (21, 21, 'neigh_op_rgt_3')
// (21, 22, 'neigh_op_bnr_3')
// (22, 19, 'local_g3_7')
// (22, 19, 'lutff_7/in_1')
// (22, 19, 'sp4_r_v_b_47')
// (22, 20, 'neigh_op_top_3')
// (22, 20, 'sp4_r_v_b_34')
// (22, 21, 'lutff_3/out')
// (22, 21, 'sp4_r_v_b_23')
// (22, 22, 'neigh_op_bot_3')
// (22, 22, 'sp4_r_v_b_10')
// (23, 18, 'sp4_v_t_47')
// (23, 19, 'sp4_v_b_47')
// (23, 20, 'neigh_op_tnl_3')
// (23, 20, 'sp4_v_b_34')
// (23, 21, 'neigh_op_lft_3')
// (23, 21, 'sp4_v_b_23')
// (23, 22, 'neigh_op_bnl_3')
// (23, 22, 'sp4_v_b_10')

reg n1694 = 0;
// (21, 20, 'sp4_r_v_b_43')
// (21, 21, 'sp4_r_v_b_30')
// (21, 22, 'neigh_op_tnr_3')
// (21, 22, 'sp4_r_v_b_19')
// (21, 23, 'neigh_op_rgt_3')
// (21, 23, 'sp4_r_v_b_6')
// (21, 24, 'neigh_op_bnr_3')
// (22, 19, 'sp4_v_t_43')
// (22, 20, 'local_g2_3')
// (22, 20, 'lutff_6/in_3')
// (22, 20, 'sp4_v_b_43')
// (22, 21, 'sp4_v_b_30')
// (22, 22, 'neigh_op_top_3')
// (22, 22, 'sp4_v_b_19')
// (22, 23, 'lutff_3/out')
// (22, 23, 'sp4_v_b_6')
// (22, 24, 'neigh_op_bot_3')
// (23, 22, 'neigh_op_tnl_3')
// (23, 23, 'neigh_op_lft_3')
// (23, 24, 'neigh_op_bnl_3')

wire n1695;
// (21, 21, 'lutff_0/lout')
// (21, 21, 'lutff_1/in_2')

wire n1696;
// (21, 21, 'lutff_1/lout')
// (21, 21, 'lutff_2/in_2')

reg n1697 = 0;
// (21, 21, 'neigh_op_tnr_1')
// (21, 22, 'neigh_op_rgt_1')
// (21, 23, 'neigh_op_bnr_1')
// (22, 19, 'sp12_v_t_22')
// (22, 20, 'sp12_v_b_22')
// (22, 21, 'neigh_op_top_1')
// (22, 21, 'sp12_v_b_21')
// (22, 22, 'lutff_1/out')
// (22, 22, 'sp12_v_b_18')
// (22, 23, 'neigh_op_bot_1')
// (22, 23, 'sp12_v_b_17')
// (22, 24, 'sp12_v_b_14')
// (22, 25, 'sp12_v_b_13')
// (22, 26, 'sp12_v_b_10')
// (22, 27, 'sp12_v_b_9')
// (22, 28, 'sp12_v_b_6')
// (22, 29, 'sp12_v_b_5')
// (22, 30, 'sp12_v_b_2')
// (22, 31, 'sp12_h_r_1')
// (22, 31, 'sp12_v_b_1')
// (23, 21, 'neigh_op_tnl_1')
// (23, 22, 'neigh_op_lft_1')
// (23, 23, 'neigh_op_bnl_1')
// (23, 31, 'sp12_h_r_2')
// (24, 31, 'sp12_h_r_5')
// (24, 31, 'sp4_h_r_2')
// (25, 31, 'sp12_h_r_6')
// (25, 31, 'sp4_h_r_15')
// (26, 31, 'sp12_h_r_9')
// (26, 31, 'sp4_h_r_26')
// (27, 31, 'sp12_h_r_10')
// (27, 31, 'sp4_h_r_39')
// (27, 32, 'sp4_r_v_b_42')
// (28, 31, 'sp12_h_r_13')
// (28, 31, 'sp4_h_l_39')
// (28, 31, 'sp4_v_t_42')
// (28, 32, 'sp4_v_b_42')
// (28, 33, 'span4_horz_r_1')
// (28, 33, 'span4_vert_31')
// (29, 31, 'sp12_h_r_14')
// (29, 33, 'span4_horz_r_5')
// (30, 31, 'sp12_h_r_17')
// (30, 33, 'span4_horz_r_9')
// (31, 31, 'sp12_h_r_18')
// (31, 33, 'io_1/D_OUT_0')
// (31, 33, 'local_g0_5')
// (31, 33, 'span4_horz_r_13')
// (32, 31, 'sp12_h_r_21')
// (32, 33, 'span4_horz_l_13')
// (33, 31, 'span12_horz_21')

reg n1698 = 0;
// (21, 21, 'sp4_r_v_b_37')
// (21, 22, 'local_g0_0')
// (21, 22, 'lutff_5/in_1')
// (21, 22, 'sp4_r_v_b_24')
// (21, 23, 'neigh_op_tnr_0')
// (21, 23, 'sp4_r_v_b_13')
// (21, 24, 'neigh_op_rgt_0')
// (21, 24, 'sp4_r_v_b_0')
// (21, 25, 'neigh_op_bnr_0')
// (22, 20, 'sp4_v_t_37')
// (22, 21, 'sp4_v_b_37')
// (22, 22, 'sp4_v_b_24')
// (22, 23, 'neigh_op_top_0')
// (22, 23, 'sp4_v_b_13')
// (22, 24, 'lutff_0/out')
// (22, 24, 'sp4_v_b_0')
// (22, 25, 'neigh_op_bot_0')
// (23, 23, 'neigh_op_tnl_0')
// (23, 24, 'neigh_op_lft_0')
// (23, 25, 'neigh_op_bnl_0')

reg n1699 = 0;
// (21, 21, 'sp4_r_v_b_44')
// (21, 22, 'local_g0_2')
// (21, 22, 'lutff_3/in_1')
// (21, 22, 'sp4_r_v_b_33')
// (21, 23, 'sp4_r_v_b_20')
// (21, 24, 'sp4_r_v_b_9')
// (22, 19, 'neigh_op_tnr_2')
// (22, 20, 'neigh_op_rgt_2')
// (22, 20, 'sp4_h_r_9')
// (22, 20, 'sp4_v_t_44')
// (22, 21, 'neigh_op_bnr_2')
// (22, 21, 'sp4_v_b_44')
// (22, 22, 'sp4_v_b_33')
// (22, 23, 'sp4_v_b_20')
// (22, 24, 'sp4_v_b_9')
// (23, 19, 'neigh_op_top_2')
// (23, 20, 'lutff_2/out')
// (23, 20, 'sp4_h_r_20')
// (23, 21, 'neigh_op_bot_2')
// (24, 19, 'neigh_op_tnl_2')
// (24, 20, 'neigh_op_lft_2')
// (24, 20, 'sp4_h_r_33')
// (24, 21, 'neigh_op_bnl_2')
// (25, 20, 'sp4_h_r_44')
// (26, 20, 'sp4_h_l_44')

reg n1700 = 0;
// (21, 22, 'local_g3_2')
// (21, 22, 'lutff_0/in_3')
// (21, 22, 'neigh_op_tnr_2')
// (21, 23, 'neigh_op_rgt_2')
// (21, 24, 'neigh_op_bnr_2')
// (22, 22, 'neigh_op_top_2')
// (22, 23, 'lutff_2/out')
// (22, 24, 'neigh_op_bot_2')
// (23, 22, 'neigh_op_tnl_2')
// (23, 23, 'neigh_op_lft_2')
// (23, 24, 'neigh_op_bnl_2')

wire n1701;
// (22, 10, 'lutff_0/cout')
// (22, 10, 'lutff_1/in_3')

wire n1702;
// (22, 10, 'lutff_1/cout')
// (22, 10, 'lutff_2/in_3')

wire n1703;
// (22, 10, 'lutff_2/cout')
// (22, 10, 'lutff_3/in_3')

wire n1704;
// (22, 10, 'lutff_3/cout')
// (22, 10, 'lutff_4/in_3')

wire n1705;
// (22, 10, 'lutff_4/cout')
// (22, 10, 'lutff_5/in_3')

wire n1706;
// (22, 10, 'lutff_5/cout')
// (22, 10, 'lutff_6/in_3')

wire n1707;
// (22, 10, 'lutff_6/cout')
// (22, 10, 'lutff_7/in_3')

wire n1708;
// (22, 10, 'lutff_7/cout')
// (22, 11, 'carry_in')
// (22, 11, 'carry_in_mux')
// (22, 11, 'lutff_0/in_3')

reg n1709 = 0;
// (22, 11, 'neigh_op_tnr_3')
// (22, 12, 'neigh_op_rgt_3')
// (22, 12, 'sp4_r_v_b_38')
// (22, 13, 'neigh_op_bnr_3')
// (22, 13, 'sp4_r_v_b_27')
// (22, 14, 'sp4_r_v_b_14')
// (22, 15, 'sp4_r_v_b_3')
// (22, 16, 'sp4_r_v_b_43')
// (22, 17, 'local_g0_6')
// (22, 17, 'lutff_1/in_1')
// (22, 17, 'sp4_r_v_b_30')
// (22, 18, 'sp4_r_v_b_19')
// (22, 19, 'sp4_r_v_b_6')
// (23, 11, 'neigh_op_top_3')
// (23, 11, 'sp4_v_t_38')
// (23, 12, 'lutff_3/out')
// (23, 12, 'sp4_v_b_38')
// (23, 13, 'neigh_op_bot_3')
// (23, 13, 'sp4_v_b_27')
// (23, 14, 'sp4_v_b_14')
// (23, 15, 'sp4_v_b_3')
// (23, 15, 'sp4_v_t_43')
// (23, 16, 'sp4_v_b_43')
// (23, 17, 'sp4_v_b_30')
// (23, 18, 'sp4_v_b_19')
// (23, 19, 'sp4_v_b_6')
// (24, 11, 'neigh_op_tnl_3')
// (24, 12, 'neigh_op_lft_3')
// (24, 13, 'neigh_op_bnl_3')

reg n1710 = 0;
// (22, 12, 'neigh_op_tnr_1')
// (22, 13, 'neigh_op_rgt_1')
// (22, 14, 'neigh_op_bnr_1')
// (23, 10, 'sp12_v_t_22')
// (23, 11, 'sp12_v_b_22')
// (23, 12, 'neigh_op_top_1')
// (23, 12, 'sp12_v_b_21')
// (23, 13, 'lutff_1/out')
// (23, 13, 'sp12_v_b_18')
// (23, 14, 'neigh_op_bot_1')
// (23, 14, 'sp12_v_b_17')
// (23, 15, 'sp12_v_b_14')
// (23, 16, 'sp12_v_b_13')
// (23, 17, 'sp12_v_b_10')
// (23, 18, 'sp12_v_b_9')
// (23, 19, 'local_g2_6')
// (23, 19, 'lutff_1/in_3')
// (23, 19, 'sp12_v_b_6')
// (23, 20, 'sp12_v_b_5')
// (23, 21, 'sp12_v_b_2')
// (23, 22, 'sp12_v_b_1')
// (24, 12, 'neigh_op_tnl_1')
// (24, 13, 'neigh_op_lft_1')
// (24, 14, 'neigh_op_bnl_1')

reg n1711 = 0;
// (22, 12, 'neigh_op_tnr_5')
// (22, 13, 'neigh_op_rgt_5')
// (22, 14, 'neigh_op_bnr_5')
// (23, 12, 'neigh_op_top_5')
// (23, 13, 'local_g2_5')
// (23, 13, 'lutff_4/in_3')
// (23, 13, 'lutff_5/out')
// (23, 14, 'neigh_op_bot_5')
// (24, 12, 'neigh_op_tnl_5')
// (24, 13, 'neigh_op_lft_5')
// (24, 14, 'neigh_op_bnl_5')

reg n1712 = 0;
// (22, 13, 'local_g1_2')
// (22, 13, 'lutff_6/in_3')
// (22, 13, 'sp4_h_r_10')
// (23, 12, 'neigh_op_tnr_1')
// (23, 13, 'neigh_op_rgt_1')
// (23, 13, 'sp4_h_r_23')
// (23, 14, 'neigh_op_bnr_1')
// (24, 12, 'neigh_op_top_1')
// (24, 13, 'lutff_1/out')
// (24, 13, 'sp4_h_r_34')
// (24, 14, 'neigh_op_bot_1')
// (25, 12, 'neigh_op_tnl_1')
// (25, 13, 'neigh_op_lft_1')
// (25, 13, 'sp4_h_r_47')
// (25, 14, 'neigh_op_bnl_1')
// (26, 13, 'sp4_h_l_47')

wire n1713;
// (22, 13, 'lutff_0/lout')
// (22, 13, 'lutff_1/in_2')

wire n1714;
// (22, 13, 'lutff_3/lout')
// (22, 13, 'lutff_4/in_2')

wire n1715;
// (22, 13, 'lutff_6/lout')
// (22, 13, 'lutff_7/in_2')

reg n1716 = 0;
// (22, 13, 'neigh_op_tnr_3')
// (22, 14, 'neigh_op_rgt_3')
// (22, 14, 'sp4_r_v_b_38')
// (22, 15, 'neigh_op_bnr_3')
// (22, 15, 'sp4_r_v_b_27')
// (22, 16, 'sp4_r_v_b_14')
// (22, 17, 'sp4_r_v_b_3')
// (23, 13, 'neigh_op_top_3')
// (23, 13, 'sp4_v_t_38')
// (23, 14, 'lutff_3/out')
// (23, 14, 'sp4_v_b_38')
// (23, 15, 'neigh_op_bot_3')
// (23, 15, 'sp4_v_b_27')
// (23, 16, 'sp4_v_b_14')
// (23, 17, 'local_g1_3')
// (23, 17, 'lutff_1/in_1')
// (23, 17, 'sp4_v_b_3')
// (24, 13, 'neigh_op_tnl_3')
// (24, 14, 'neigh_op_lft_3')
// (24, 15, 'neigh_op_bnl_3')

reg n1717 = 0;
// (22, 13, 'neigh_op_tnr_4')
// (22, 14, 'neigh_op_rgt_4')
// (22, 14, 'sp4_r_v_b_40')
// (22, 15, 'neigh_op_bnr_4')
// (22, 15, 'sp4_r_v_b_29')
// (22, 16, 'sp4_r_v_b_16')
// (22, 17, 'sp4_r_v_b_5')
// (23, 13, 'neigh_op_top_4')
// (23, 13, 'sp4_v_t_40')
// (23, 14, 'lutff_4/out')
// (23, 14, 'sp4_v_b_40')
// (23, 15, 'neigh_op_bot_4')
// (23, 15, 'sp4_v_b_29')
// (23, 16, 'sp4_v_b_16')
// (23, 17, 'local_g1_5')
// (23, 17, 'lutff_3/in_1')
// (23, 17, 'sp4_v_b_5')
// (24, 13, 'neigh_op_tnl_4')
// (24, 14, 'neigh_op_lft_4')
// (24, 15, 'neigh_op_bnl_4')

reg n1718 = 0;
// (22, 13, 'neigh_op_tnr_5')
// (22, 14, 'neigh_op_rgt_5')
// (22, 14, 'sp4_r_v_b_42')
// (22, 15, 'neigh_op_bnr_5')
// (22, 15, 'sp4_r_v_b_31')
// (22, 16, 'sp4_r_v_b_18')
// (22, 17, 'sp4_r_v_b_7')
// (23, 13, 'neigh_op_top_5')
// (23, 13, 'sp4_v_t_42')
// (23, 14, 'lutff_5/out')
// (23, 14, 'sp4_v_b_42')
// (23, 15, 'neigh_op_bot_5')
// (23, 15, 'sp4_v_b_31')
// (23, 16, 'sp4_v_b_18')
// (23, 17, 'local_g0_7')
// (23, 17, 'lutff_6/in_1')
// (23, 17, 'sp4_v_b_7')
// (24, 13, 'neigh_op_tnl_5')
// (24, 14, 'neigh_op_lft_5')
// (24, 15, 'neigh_op_bnl_5')

reg n1719 = 0;
// (22, 14, 'neigh_op_tnr_3')
// (22, 15, 'neigh_op_rgt_3')
// (22, 15, 'sp4_r_v_b_38')
// (22, 16, 'neigh_op_bnr_3')
// (22, 16, 'sp4_r_v_b_27')
// (22, 17, 'sp4_r_v_b_14')
// (22, 18, 'sp4_r_v_b_3')
// (23, 14, 'neigh_op_top_3')
// (23, 14, 'sp4_v_t_38')
// (23, 15, 'lutff_3/out')
// (23, 15, 'sp4_v_b_38')
// (23, 16, 'neigh_op_bot_3')
// (23, 16, 'sp4_v_b_27')
// (23, 17, 'local_g0_6')
// (23, 17, 'lutff_1/in_3')
// (23, 17, 'sp4_v_b_14')
// (23, 18, 'sp4_v_b_3')
// (24, 14, 'neigh_op_tnl_3')
// (24, 15, 'neigh_op_lft_3')
// (24, 16, 'neigh_op_bnl_3')

reg n1720 = 0;
// (22, 14, 'neigh_op_tnr_4')
// (22, 15, 'neigh_op_rgt_4')
// (22, 16, 'neigh_op_bnr_4')
// (23, 14, 'neigh_op_top_4')
// (23, 15, 'lutff_4/out')
// (23, 15, 'sp4_r_v_b_41')
// (23, 16, 'neigh_op_bot_4')
// (23, 16, 'sp4_r_v_b_28')
// (23, 17, 'local_g3_1')
// (23, 17, 'lutff_3/in_3')
// (23, 17, 'sp4_r_v_b_17')
// (23, 18, 'sp4_r_v_b_4')
// (24, 14, 'neigh_op_tnl_4')
// (24, 14, 'sp4_v_t_41')
// (24, 15, 'neigh_op_lft_4')
// (24, 15, 'sp4_v_b_41')
// (24, 16, 'neigh_op_bnl_4')
// (24, 16, 'sp4_v_b_28')
// (24, 17, 'sp4_v_b_17')
// (24, 18, 'sp4_v_b_4')

reg n1721 = 0;
// (22, 14, 'neigh_op_tnr_5')
// (22, 15, 'neigh_op_rgt_5')
// (22, 15, 'sp4_r_v_b_42')
// (22, 16, 'neigh_op_bnr_5')
// (22, 16, 'sp4_r_v_b_31')
// (22, 17, 'sp4_r_v_b_18')
// (22, 18, 'sp4_r_v_b_7')
// (23, 14, 'neigh_op_top_5')
// (23, 14, 'sp4_v_t_42')
// (23, 15, 'lutff_5/out')
// (23, 15, 'sp4_v_b_42')
// (23, 16, 'neigh_op_bot_5')
// (23, 16, 'sp4_v_b_31')
// (23, 17, 'local_g1_2')
// (23, 17, 'lutff_6/in_3')
// (23, 17, 'sp4_v_b_18')
// (23, 18, 'sp4_v_b_7')
// (24, 14, 'neigh_op_tnl_5')
// (24, 15, 'neigh_op_lft_5')
// (24, 16, 'neigh_op_bnl_5')

wire n1722;
// (22, 16, 'lutff_1/lout')
// (22, 16, 'lutff_2/in_2')

wire n1723;
// (22, 16, 'lutff_3/lout')
// (22, 16, 'lutff_4/in_2')

wire n1724;
// (22, 16, 'lutff_5/lout')
// (22, 16, 'lutff_6/in_2')

wire n1725;
// (22, 16, 'lutff_6/lout')
// (22, 16, 'lutff_7/in_2')

reg n1726 = 0;
// (22, 16, 'neigh_op_tnr_0')
// (22, 17, 'neigh_op_rgt_0')
// (22, 18, 'neigh_op_bnr_0')
// (23, 16, 'neigh_op_top_0')
// (23, 17, 'local_g1_0')
// (23, 17, 'lutff_0/out')
// (23, 17, 'lutff_2/in_3')
// (23, 18, 'neigh_op_bot_0')
// (24, 16, 'neigh_op_tnl_0')
// (24, 17, 'neigh_op_lft_0')
// (24, 18, 'neigh_op_bnl_0')

wire n1727;
// (22, 16, 'neigh_op_tnr_2')
// (22, 17, 'local_g3_2')
// (22, 17, 'lutff_4/in_3')
// (22, 17, 'neigh_op_rgt_2')
// (22, 18, 'neigh_op_bnr_2')
// (23, 16, 'neigh_op_top_2')
// (23, 17, 'lutff_2/out')
// (23, 18, 'neigh_op_bot_2')
// (24, 16, 'neigh_op_tnl_2')
// (24, 17, 'neigh_op_lft_2')
// (24, 18, 'neigh_op_bnl_2')

wire n1728;
// (22, 16, 'neigh_op_tnr_4')
// (22, 17, 'neigh_op_rgt_4')
// (22, 18, 'local_g0_4')
// (22, 18, 'lutff_3/in_3')
// (22, 18, 'neigh_op_bnr_4')
// (23, 16, 'neigh_op_top_4')
// (23, 17, 'lutff_4/out')
// (23, 18, 'neigh_op_bot_4')
// (24, 16, 'neigh_op_tnl_4')
// (24, 17, 'neigh_op_lft_4')
// (24, 18, 'neigh_op_bnl_4')

reg n1729 = 0;
// (22, 16, 'neigh_op_tnr_5')
// (22, 17, 'neigh_op_rgt_5')
// (22, 18, 'neigh_op_bnr_5')
// (23, 16, 'neigh_op_top_5')
// (23, 17, 'local_g2_5')
// (23, 17, 'lutff_4/in_3')
// (23, 17, 'lutff_5/out')
// (23, 18, 'neigh_op_bot_5')
// (24, 16, 'neigh_op_tnl_5')
// (24, 17, 'neigh_op_lft_5')
// (24, 18, 'neigh_op_bnl_5')

wire n1730;
// (22, 17, 'lutff_0/lout')
// (22, 17, 'lutff_1/in_2')

wire n1731;
// (22, 17, 'lutff_2/lout')
// (22, 17, 'lutff_3/in_2')

wire n1732;
// (22, 17, 'lutff_4/lout')
// (22, 17, 'lutff_5/in_2')

reg n1733 = 0;
// (22, 17, 'neigh_op_tnr_0')
// (22, 18, 'neigh_op_rgt_0')
// (22, 19, 'local_g1_0')
// (22, 19, 'lutff_6/in_3')
// (22, 19, 'neigh_op_bnr_0')
// (23, 17, 'neigh_op_top_0')
// (23, 18, 'lutff_0/out')
// (23, 19, 'neigh_op_bot_0')
// (24, 17, 'neigh_op_tnl_0')
// (24, 18, 'neigh_op_lft_0')
// (24, 19, 'neigh_op_bnl_0')

reg n1734 = 0;
// (22, 17, 'neigh_op_tnr_2')
// (22, 18, 'neigh_op_rgt_2')
// (22, 19, 'local_g0_2')
// (22, 19, 'lutff_7/in_3')
// (22, 19, 'neigh_op_bnr_2')
// (23, 17, 'neigh_op_top_2')
// (23, 18, 'lutff_2/out')
// (23, 19, 'neigh_op_bot_2')
// (24, 17, 'neigh_op_tnl_2')
// (24, 18, 'neigh_op_lft_2')
// (24, 19, 'neigh_op_bnl_2')

wire n1735;
// (22, 17, 'sp4_r_v_b_42')
// (22, 18, 'local_g0_7')
// (22, 18, 'lutff_4/in_1')
// (22, 18, 'neigh_op_tnr_1')
// (22, 18, 'sp4_r_v_b_31')
// (22, 19, 'neigh_op_rgt_1')
// (22, 19, 'sp4_r_v_b_18')
// (22, 20, 'neigh_op_bnr_1')
// (22, 20, 'sp4_r_v_b_7')
// (23, 16, 'sp4_v_t_42')
// (23, 17, 'sp4_v_b_42')
// (23, 18, 'neigh_op_top_1')
// (23, 18, 'sp4_v_b_31')
// (23, 19, 'lutff_1/out')
// (23, 19, 'sp4_v_b_18')
// (23, 20, 'neigh_op_bot_1')
// (23, 20, 'sp4_v_b_7')
// (24, 18, 'neigh_op_tnl_1')
// (24, 19, 'neigh_op_lft_1')
// (24, 20, 'neigh_op_bnl_1')

wire n1736;
// (22, 18, 'lutff_0/lout')
// (22, 18, 'lutff_1/in_2')

wire n1737;
// (22, 18, 'lutff_1/lout')
// (22, 18, 'lutff_2/in_2')

wire n1738;
// (22, 18, 'lutff_4/lout')
// (22, 18, 'lutff_5/in_2')

wire n1739;
// (22, 18, 'lutff_5/lout')
// (22, 18, 'lutff_6/in_2')

wire n1740;
// (22, 20, 'lutff_2/lout')
// (22, 20, 'lutff_3/in_2')

wire n1741;
// (22, 20, 'lutff_3/lout')
// (22, 20, 'lutff_4/in_2')

reg n1742 = 0;
// (23, 13, 'local_g3_0')
// (23, 13, 'lutff_4/in_1')
// (23, 13, 'sp4_r_v_b_40')
// (23, 14, 'sp4_r_v_b_29')
// (23, 15, 'sp4_r_v_b_16')
// (23, 16, 'neigh_op_tnr_6')
// (23, 16, 'sp4_r_v_b_5')
// (23, 17, 'neigh_op_rgt_6')
// (23, 17, 'sp4_r_v_b_44')
// (23, 18, 'neigh_op_bnr_6')
// (23, 18, 'sp4_r_v_b_33')
// (23, 19, 'sp4_r_v_b_20')
// (23, 20, 'sp4_r_v_b_9')
// (24, 12, 'sp4_v_t_40')
// (24, 13, 'sp4_v_b_40')
// (24, 14, 'sp4_v_b_29')
// (24, 15, 'sp4_v_b_16')
// (24, 16, 'neigh_op_top_6')
// (24, 16, 'sp4_v_b_5')
// (24, 16, 'sp4_v_t_44')
// (24, 17, 'lutff_6/out')
// (24, 17, 'sp4_v_b_44')
// (24, 18, 'neigh_op_bot_6')
// (24, 18, 'sp4_v_b_33')
// (24, 19, 'sp4_v_b_20')
// (24, 20, 'sp4_v_b_9')
// (25, 16, 'neigh_op_tnl_6')
// (25, 17, 'neigh_op_lft_6')
// (25, 18, 'neigh_op_bnl_6')

reg n1743 = 0;
// (23, 15, 'neigh_op_tnr_1')
// (23, 16, 'neigh_op_rgt_1')
// (23, 17, 'local_g1_1')
// (23, 17, 'lutff_7/in_3')
// (23, 17, 'neigh_op_bnr_1')
// (24, 15, 'neigh_op_top_1')
// (24, 16, 'lutff_1/out')
// (24, 17, 'neigh_op_bot_1')
// (25, 15, 'neigh_op_tnl_1')
// (25, 16, 'neigh_op_lft_1')
// (25, 17, 'neigh_op_bnl_1')

reg n1744 = 0;
// (23, 16, 'neigh_op_tnr_4')
// (23, 17, 'neigh_op_rgt_4')
// (23, 17, 'sp4_r_v_b_40')
// (23, 18, 'neigh_op_bnr_4')
// (23, 18, 'sp4_r_v_b_29')
// (23, 19, 'local_g3_0')
// (23, 19, 'lutff_1/in_0')
// (23, 19, 'sp4_r_v_b_16')
// (23, 20, 'sp4_r_v_b_5')
// (24, 16, 'neigh_op_top_4')
// (24, 16, 'sp4_v_t_40')
// (24, 17, 'lutff_4/out')
// (24, 17, 'sp4_v_b_40')
// (24, 18, 'neigh_op_bot_4')
// (24, 18, 'sp4_v_b_29')
// (24, 19, 'sp4_v_b_16')
// (24, 20, 'sp4_v_b_5')
// (25, 16, 'neigh_op_tnl_4')
// (25, 17, 'neigh_op_lft_4')
// (25, 18, 'neigh_op_bnl_4')

wire n1745;
// (23, 17, 'lutff_1/lout')
// (23, 17, 'lutff_2/in_2')

wire n1746;
// (23, 17, 'lutff_3/lout')
// (23, 17, 'lutff_4/in_2')

wire n1747;
// (23, 17, 'lutff_6/lout')
// (23, 17, 'lutff_7/in_2')

wire io_33_27_1;
// (23, 21, 'neigh_op_tnr_4')
// (23, 22, 'neigh_op_rgt_4')
// (23, 23, 'neigh_op_bnr_4')
// (24, 21, 'neigh_op_top_4')
// (24, 22, 'lutff_4/out')
// (24, 22, 'sp4_r_v_b_41')
// (24, 23, 'neigh_op_bot_4')
// (24, 23, 'sp4_r_v_b_28')
// (24, 24, 'sp4_r_v_b_17')
// (24, 25, 'sp4_r_v_b_4')
// (25, 21, 'neigh_op_tnl_4')
// (25, 21, 'sp4_v_t_41')
// (25, 22, 'neigh_op_lft_4')
// (25, 22, 'sp4_v_b_41')
// (25, 23, 'neigh_op_bnl_4')
// (25, 23, 'sp4_v_b_28')
// (25, 24, 'sp4_v_b_17')
// (25, 25, 'sp4_h_r_10')
// (25, 25, 'sp4_v_b_4')
// (26, 25, 'sp4_h_r_23')
// (27, 25, 'sp4_h_r_34')
// (28, 25, 'sp4_h_r_47')
// (29, 25, 'sp4_h_l_47')
// (29, 25, 'sp4_h_r_6')
// (30, 25, 'sp4_h_r_19')
// (31, 25, 'sp4_h_r_30')
// (32, 25, 'sp4_h_r_43')
// (33, 25, 'span4_horz_43')
// (33, 25, 'span4_vert_t_15')
// (33, 26, 'span4_vert_b_15')
// (33, 27, 'io_1/D_OUT_0')
// (33, 27, 'io_1/PAD')
// (33, 27, 'local_g0_3')
// (33, 27, 'span4_vert_b_11')
// (33, 28, 'span4_vert_b_7')
// (33, 29, 'span4_vert_b_3')

wire io_26_33_1;
// (26, 33, 'io_1/D_OUT_0')
// (26, 33, 'io_1/PAD')

wire io_27_33_0;
// (27, 33, 'io_0/PAD')

wire io_28_33_1;
// (28, 33, 'io_1/PAD')

wire io_29_33_0;
// (29, 33, 'io_0/PAD')

wire io_29_33_1;
// (29, 33, 'io_1/PAD')

wire io_30_0_0;
// (30, 0, 'io_0/D_OUT_0')
// (30, 0, 'io_0/PAD')

wire io_30_33_0;
// (30, 33, 'io_0/PAD')

wire io_30_33_1;
// (30, 33, 'io_1/PAD')

wire io_31_0_0;
// (31, 0, 'io_0/D_OUT_0')
// (31, 0, 'io_0/PAD')

wire io_31_0_1;
// (31, 0, 'io_1/D_OUT_0')
// (31, 0, 'io_1/PAD')

wire io_31_33_0;
// (31, 33, 'io_0/PAD')

wire io_31_33_1;
// (31, 33, 'io_1/PAD')

wire io_33_2_1;
// (33, 2, 'io_1/PAD')

wire io_33_6_1;
// (33, 6, 'io_1/PAD')

wire io_33_10_1;
// (33, 10, 'io_1/PAD')

wire io_33_14_1;
// (33, 14, 'io_1/PAD')

wire io_33_15_0;
// (33, 15, 'io_0/PAD')

wire io_33_15_1;
// (33, 15, 'io_1/PAD')

wire io_33_16_0;
// (33, 16, 'io_0/PAD')

wire io_33_16_1;
// (33, 16, 'io_1/PAD')

wire io_33_17_0;
// (33, 17, 'io_0/D_OUT_0')
// (33, 17, 'io_0/PAD')

wire io_33_19_1;
// (33, 19, 'io_1/D_OUT_0')
// (33, 19, 'io_1/PAD')

wire io_33_20_1;
// (33, 20, 'io_1/D_OUT_0')
// (33, 20, 'io_1/PAD')

wire n1772;
// (1, 1, 'neigh_op_bnl_1')

wire n1773;
// (32, 1, 'neigh_op_bnr_3')

wire n1774;
// (17, 20, 'lutff_6/cout')

wire n1775;
// (12, 22, 'lutff_5/cout')

wire n1776;
// (11, 20, 'lutff_1/cout')

wire n1777;
// (17, 24, 'lutff_6/cout')

wire n1778;
// (12, 21, 'lutff_4/cout')

wire n1779;
// (17, 22, 'lutff_4/cout')

wire n1780;
// (12, 15, 'lutff_2/cout')

wire n1781;
// (15, 21, 'lutff_4/cout')

wire n1782;
// (15, 22, 'lutff_6/cout')

wire n1783;
// (17, 23, 'lutff_3/cout')

wire n1784;
// (12, 14, 'lutff_1/cout')

wire n1785;
// (11, 19, 'lutff_4/cout')

wire n1786;
// (13, 18, 'lutff_3/cout')

wire n1787;
// (15, 20, 'lutff_4/cout')

wire n1788;
// (13, 19, 'lutff_4/cout')

wire n1789;
// (17, 18, 'lutff_0/cout')

wire n1790;
// (13, 23, 'lutff_1/cout')

wire n1791;
// (13, 20, 'lutff_5/cout')

wire n1792;
// (13, 24, 'lutff_0/cout')

wire n1793;
// (11, 20, 'lutff_4/cout')

wire n1794;
// (11, 18, 'lutff_2/cout')

wire n1795;
// (17, 20, 'lutff_2/cout')

wire n1796;
// (11, 19, 'lutff_1/cout')

wire n1797;
// (13, 18, 'lutff_6/cout')

wire n1798;
// (17, 22, 'lutff_0/cout')

wire n1799;
// (12, 15, 'lutff_6/cout')

wire n1800;
// (13, 19, 'lutff_1/cout')

wire n1801;
// (15, 21, 'lutff_0/cout')

wire n1802;
// (13, 23, 'lutff_6/cout')

wire n1803;
// (12, 14, 'lutff_5/cout')

wire n1804;
// (10, 10, 'lutff_4/cout')

wire n1805;
// (10, 17, 'lutff_6/cout')

wire n1806;
// (13, 20, 'lutff_0/cout')

wire n1807;
// (17, 19, 'lutff_4/cout')

wire n1808;
// (13, 22, 'lutff_2/cout')

wire n1809;
// (17, 18, 'lutff_4/cout')

wire n1810;
// (12, 23, 'lutff_1/cout')

wire n1811;
// (12, 22, 'lutff_2/cout')

wire n1812;
// (11, 20, 'lutff_0/cout')

wire n1813;
// (17, 24, 'lutff_1/cout')

wire n1814;
// (12, 21, 'lutff_3/cout')

wire n1815;
// (15, 21, 'lutff_5/cout')

wire n1816;
// (11, 18, 'lutff_6/cout')

wire n1817;
// (15, 22, 'lutff_1/cout')

wire n1818;
// (11, 19, 'lutff_5/cout')

wire n1819;
// (13, 18, 'lutff_2/cout')

wire n1820;
// (15, 20, 'lutff_3/cout')

wire n1821;
// (13, 19, 'lutff_5/cout')

wire n1822;
// (13, 23, 'lutff_2/cout')

wire n1823;
// (13, 20, 'lutff_4/cout')

wire n1824;
// (17, 19, 'lutff_0/cout')

wire n1825;
// (13, 24, 'lutff_3/cout')

wire n1826;
// (13, 22, 'lutff_6/cout')

wire n1827;
// (12, 23, 'lutff_5/cout')

wire n1828;
// (17, 20, 'lutff_5/cout')

wire n1829;
// (12, 22, 'lutff_6/cout')

wire n1830;
// (17, 24, 'lutff_5/cout')

wire n1831;
// (13, 18, 'lutff_5/cout')

wire n1832;
// (12, 15, 'lutff_1/cout')

wire n1833;
// (13, 19, 'lutff_2/cout')

wire n1834;
// (15, 21, 'lutff_1/cout')

wire n1835;
// (15, 22, 'lutff_5/cout')

wire n1836;
// (17, 23, 'lutff_0/cout')

wire n1837;
// (12, 14, 'lutff_2/cout')

wire n1838;
// (10, 10, 'lutff_5/cout')

wire n1839;
// (13, 20, 'lutff_3/cout')

wire n1840;
// (17, 19, 'lutff_5/cout')

wire n1841;
// (13, 24, 'lutff_6/cout')

wire n1842;
// (13, 22, 'lutff_1/cout')

wire n1843;
// (17, 18, 'lutff_3/cout')

wire n1844;
// (12, 23, 'lutff_0/cout')

wire n1845;
// (12, 22, 'lutff_3/cout')

wire n1846;
// (17, 24, 'lutff_0/cout')

wire n1847;
// (12, 21, 'lutff_2/cout')

wire n1848;
// (15, 21, 'lutff_6/cout')

wire n1849;
// (11, 18, 'lutff_1/cout')

wire n1850;
// (15, 22, 'lutff_0/cout')

wire n1851;
// (17, 20, 'lutff_1/cout')

wire n1852;
// (11, 19, 'lutff_2/cout')

wire n1853;
// (13, 18, 'lutff_1/cout')

wire n1854;
// (15, 20, 'lutff_2/cout')

wire n1855;
// (17, 22, 'lutff_3/cout')

wire n1856;
// (12, 15, 'lutff_5/cout')

wire n1857;
// (13, 19, 'lutff_6/cout')

wire n1858;
// (17, 23, 'lutff_4/cout')

wire n1859;
// (13, 23, 'lutff_3/cout')

wire n1860;
// (12, 14, 'lutff_6/cout')

wire n1861;
// (10, 17, 'lutff_5/cout')

wire n1862;
// (17, 19, 'lutff_1/cout')

wire n1863;
// (13, 24, 'lutff_2/cout')

wire n1864;
// (13, 22, 'lutff_5/cout')

wire n1865;
// (12, 23, 'lutff_4/cout')

wire n1866;
// (17, 20, 'lutff_4/cout')

wire n1867;
// (11, 20, 'lutff_3/cout')

wire n1868;
// (17, 24, 'lutff_4/cout')

wire n1869;
// (12, 21, 'lutff_6/cout')

wire n1870;
// (13, 18, 'lutff_4/cout')

wire n1871;
// (17, 22, 'lutff_6/cout')

wire n1872;
// (12, 15, 'lutff_0/cout')

wire n1873;
// (13, 19, 'lutff_3/cout')

wire n1874;
// (15, 21, 'lutff_2/cout')

wire n1875;
// (11, 18, 'lutff_5/cout')

wire n1876;
// (15, 22, 'lutff_4/cout')

wire n1877;
// (17, 23, 'lutff_1/cout')

wire n1878;
// (12, 14, 'lutff_3/cout')

wire n1879;
// (10, 10, 'lutff_6/cout')

wire n1880;
// (13, 20, 'lutff_2/cout')

wire n1881;
// (17, 19, 'lutff_6/cout')

wire n1882;
// (11, 19, 'lutff_6/cout')

wire n1883;
// (15, 20, 'lutff_6/cout')

wire n1884;
// (13, 22, 'lutff_0/cout')

wire n1885;
// (17, 18, 'lutff_2/cout')

wire n1886;
// (12, 23, 'lutff_3/cout')

wire n1887;
// (12, 22, 'lutff_0/cout')

wire n1888;
// (11, 20, 'lutff_6/cout')

wire n1889;
// (17, 24, 'lutff_3/cout')

wire n1890;
// (12, 21, 'lutff_1/cout')

wire n1891;
// (11, 18, 'lutff_0/cout')

wire n1892;
// (15, 22, 'lutff_3/cout')

wire n1893;
// (17, 20, 'lutff_0/cout')

wire n1894;
// (11, 19, 'lutff_3/cout')

wire n1895;
// (13, 18, 'lutff_0/cout')

wire n1896;
// (15, 20, 'lutff_1/cout')

wire n1897;
// (17, 22, 'lutff_2/cout')

wire n1898;
// (12, 15, 'lutff_4/cout')

wire n1899;
// (17, 23, 'lutff_5/cout')

wire n1900;
// (13, 23, 'lutff_4/cout')

wire n1901;
// (13, 20, 'lutff_6/cout')

wire n1902;
// (17, 19, 'lutff_2/cout')

wire n1903;
// (13, 24, 'lutff_5/cout')

wire n1904;
// (13, 22, 'lutff_4/cout')

wire n1905;
// (17, 18, 'lutff_6/cout')

wire n1906;
// (12, 22, 'lutff_4/cout')

wire n1907;
// (11, 20, 'lutff_2/cout')

wire n1908;
// (12, 21, 'lutff_5/cout')

wire n1909;
// (17, 22, 'lutff_5/cout')

wire n1910;
// (12, 15, 'lutff_3/cout')

wire n1911;
// (15, 21, 'lutff_3/cout')

wire n1912;
// (11, 18, 'lutff_4/cout')

wire n1913;
// (17, 23, 'lutff_2/cout')

wire n1914;
// (12, 14, 'lutff_0/cout')

wire n1915;
// (15, 20, 'lutff_5/cout')

wire n1916;
// (17, 18, 'lutff_1/cout')

wire n1917;
// (13, 23, 'lutff_0/cout')

wire n1918;
// (12, 23, 'lutff_2/cout')

wire n1919;
// (13, 24, 'lutff_1/cout')

wire n1920;
// (12, 22, 'lutff_1/cout')

wire n1921;
// (11, 20, 'lutff_5/cout')

wire n1922;
// (17, 24, 'lutff_2/cout')

wire n1923;
// (12, 21, 'lutff_0/cout')

wire n1924;
// (11, 18, 'lutff_3/cout')

wire n1925;
// (15, 22, 'lutff_2/cout')

wire n1926;
// (17, 20, 'lutff_3/cout')

wire n1927;
// (11, 19, 'lutff_0/cout')

wire n1928;
// (15, 20, 'lutff_0/cout')

wire n1929;
// (17, 22, 'lutff_1/cout')

wire n1930;
// (13, 19, 'lutff_0/cout')

wire n1931;
// (17, 23, 'lutff_6/cout')

wire n1932;
// (13, 23, 'lutff_5/cout')

wire n1933;
// (12, 14, 'lutff_4/cout')

wire n1934;
// (13, 20, 'lutff_1/cout')

wire n1935;
// (17, 19, 'lutff_3/cout')

wire n1936;
// (13, 24, 'lutff_4/cout')

wire n1937;
// (13, 22, 'lutff_3/cout')

wire n1938;
// (17, 18, 'lutff_5/cout')

wire n1939;
// (12, 23, 'lutff_6/cout')

wire n1940;
// (16, 16, 'lutff_2/lout')

wire n1941;
// (22, 12, 'lutff_4/lout')

wire n1942;
// (15, 13, 'lutff_0/out')

wire n1943;
// (20, 20, 'lutff_3/lout')

wire n1944;
// (16, 14, 'lutff_7/lout')

wire n1945;
// (5, 17, 'lutff_5/lout')

wire n1946;
// (16, 19, 'lutff_4/lout')

wire n1947;
// (15, 19, 'lutff_1/lout')

wire n1948;
// (17, 20, 'lutff_6/lout')

wire n1949;
// (23, 15, 'lutff_1/lout')

wire n1950;
// (24, 16, 'lutff_1/lout')

wire n1951;
// (7, 16, 'lutff_7/lout')

wire n1952;
// (21, 11, 'lutff_0/lout')

wire n1953;
// (12, 22, 'lutff_5/out')

wire n1954;
// (12, 22, 'lutff_5/lout')

wire n1955;
// (19, 23, 'lutff_3/lout')

wire n1956;
// (10, 9, 'lutff_5/lout')

wire n1957;
// (22, 15, 'lutff_5/lout')

wire n1958;
// (20, 11, 'lutff_2/lout')

wire n1959;
// (19, 24, 'lutff_7/lout')

wire n1960;
// (11, 20, 'lutff_1/lout')

wire n1961;
// (5, 18, 'lutff_4/lout')

wire n1962;
// (16, 18, 'lutff_7/lout')

wire n1963;
// (10, 20, 'lutff_0/lout')

wire n1964;
// (21, 15, 'lutff_5/lout')

wire n1965;
// (20, 22, 'lutff_4/lout')

wire n1966;
// (17, 21, 'lutff_5/lout')

wire n1967;
// (17, 24, 'lutff_6/out')

wire n1968;
// (17, 24, 'lutff_6/lout')

wire n1969;
// (23, 12, 'lutff_0/lout')

wire n1970;
// (24, 15, 'lutff_0/lout')

wire n1971;
// (21, 12, 'lutff_1/lout')

wire n1972;
// (12, 21, 'lutff_4/lout')

wire n1973;
// (17, 10, 'lutff_1/lout')

wire n1974;
// (19, 20, 'lutff_2/lout')

wire n1975;
// (22, 14, 'lutff_2/lout')

wire n1976;
// (23, 16, 'lutff_6/lout')

wire n1977;
// (11, 14, 'lutff_7/lout')

wire n1978;
// (16, 12, 'lutff_1/lout')

wire n1979;
// (16, 17, 'lutff_6/lout')

wire n1980;
// (13, 15, 'lutff_0/lout')

wire n1981;
// (15, 17, 'lutff_7/lout')

wire n1982;
// (20, 24, 'lutff_2/lout')

wire n1983;
// (20, 21, 'lutff_5/lout')

wire n1984;
// (17, 22, 'lutff_4/lout')

wire n1985;
// (24, 14, 'lutff_3/lout')

wire n1986;
// (22, 10, 'lutff_7/lout')

wire n1987;
// (21, 13, 'lutff_2/out')

wire n1988;
// (12, 15, 'lutff_2/lout')

wire n1989;
// (19, 21, 'lutff_5/lout')

wire n1990;
// (16, 8, 'lutff_6/lout')

wire n1991;
// (24, 17, 'lutff_7/lout')

wire n1992;
// (15, 21, 'lutff_4/lout')

wire n1993;
// (23, 17, 'lutff_1/out')

wire n1994;
// (11, 15, 'lutff_4/lout')

wire n1995;
// (11, 18, 'lutff_7/lout')

wire n1996;
// (16, 11, 'lutff_0/lout')

wire n1997;
// (13, 16, 'lutff_1/lout')

wire n1998;
// (15, 22, 'lutff_6/out')

wire n1999;
// (15, 22, 'lutff_6/lout')

wire n2000;
// (18, 9, 'lutff_2/lout')

wire n2001;
// (6, 11, 'lutff_5/lout')

wire n2002;
// (12, 24, 'lutff_0/lout')

wire n2003;
// (17, 23, 'lutff_3/lout')

wire n2004;
// (19, 17, 'lutff_2/lout')

wire n2005;
// (22, 21, 'lutff_5/lout')

wire n2006;
// (24, 13, 'lutff_2/lout')

wire n2007;
// (21, 14, 'lutff_3/out')

wire n2008;
// (9, 16, 'lutff_0/lout')

wire n2009;
// (12, 14, 'lutff_1/lout')

wire n2010;
// (14, 20, 'lutff_0/lout')

wire n2011;
// (19, 18, 'lutff_4/out')

wire n2012;
// (10, 10, 'lutff_0/out')

wire n2013;
// (10, 10, 'lutff_0/lout')

wire n2014;
// (10, 10, 'carry_in_mux')

// Carry-In for (10 10)
assign n2014 = 0;

wire n2015;
// (16, 23, 'lutff_7/lout')

wire n2016;
// (15, 10, 'lutff_5/lout')

wire n2017;
// (20, 19, 'lutff_6/lout')

wire n2018;
// (18, 22, 'lutff_0/lout')

wire n2019;
// (11, 12, 'lutff_5/lout')

wire n2020;
// (11, 19, 'lutff_4/lout')

wire n2021;
// (16, 10, 'lutff_3/lout')

wire n2022;
// (9, 12, 'lutff_2/out')

wire n2023;
// (15, 24, 'lutff_4/lout')

wire n2024;
// (13, 17, 'lutff_2/out')

wire n2025;
// (17, 16, 'lutff_2/out')

wire n2026;
// (19, 14, 'lutff_3/out')

wire n2027;
// (22, 20, 'lutff_6/lout')

wire n2028;
// (16, 24, 'lutff_3/lout')

wire n2029;
// (12, 13, 'lutff_0/lout')

wire n2030;
// (20, 12, 'lutff_4/lout')

wire n2031;
// (10, 13, 'lutff_1/lout')

wire n2032;
// (16, 22, 'lutff_4/lout')

wire n2033;
// (15, 11, 'lutff_6/lout')

wire n2034;
// (20, 18, 'lutff_5/lout')

wire n2035;
// (20, 15, 'lutff_6/lout')

wire n2036;
// (11, 13, 'lutff_2/lout')

wire n2037;
// (11, 16, 'lutff_5/lout')

wire n2038;
// (9, 13, 'lutff_1/lout')

wire n2039;
// (15, 25, 'lutff_3/lout')

wire n2040;
// (13, 18, 'lutff_3/lout')

wire n2041;
// (18, 11, 'lutff_0/lout')

wire n2042;
// (15, 20, 'lutff_4/lout')

wire n2043;
// (17, 17, 'lutff_1/out')

wire n2044;
// (16, 7, 'lutff_1/lout')

wire n2045;
// (19, 15, 'lutff_0/lout')

wire n2046;
// (22, 23, 'lutff_7/lout')

wire n2047;
// (9, 18, 'lutff_2/lout')

wire n2048;
// (11, 9, 'lutff_7/lout')

wire n2049;
// (19, 16, 'lutff_6/lout')

wire n2050;
// (16, 21, 'lutff_5/lout')

wire n2051;
// (15, 8, 'lutff_7/lout')

wire n2052;
// (6, 12, 'lutff_5/lout')

wire n2053;
// (15, 7, 'lutff_6/lout')

wire n2054;
// (18, 24, 'lutff_2/lout')

wire n2055;
// (20, 17, 'lutff_4/lout')

wire n2056;
// (20, 14, 'lutff_5/lout')

wire n2057;
// (23, 20, 'lutff_2/lout')

wire n2058;
// (11, 10, 'lutff_3/lout')

wire n2059;
// (13, 19, 'lutff_4/lout')

wire n2060;
// (14, 18, 'lutff_3/lout')

wire n2061;
// (17, 18, 'lutff_0/out')

wire n2062;
// (17, 18, 'lutff_0/lout')

wire n2063;
// (17, 18, 'carry_in_mux')

// Carry-In for (17 18)
assign n2063 = 0;

wire n2064;
// (19, 12, 'lutff_1/lout')

wire n2065;
// (17, 12, 'lutff_3/lout')

wire n2066;
// (10, 15, 'lutff_3/lout')

wire n2067;
// (16, 20, 'lutff_2/lout')

wire n2068;
// (13, 23, 'lutff_1/out')

wire n2069;
// (13, 23, 'lutff_1/lout')

wire n2070;
// (15, 9, 'lutff_0/lout')

wire n2071;
// (18, 14, 'lutff_4/out')

wire n2072;
// (20, 16, 'lutff_3/lout')

wire n2073;
// (20, 13, 'lutff_4/lout')

wire n2074;
// (11, 11, 'lutff_0/lout')

// Carry-In for (11 11)
assign n415 = 1;

wire n2075;
// (22, 18, 'lutff_5/out')

wire n2076;
// (10, 17, 'lutff_3/lout')

wire n2077;
// (9, 15, 'lutff_7/lout')

wire n2078;
// (13, 20, 'lutff_5/lout')

wire n2079;
// (18, 13, 'lutff_6/out')

wire n2080;
// (14, 13, 'lutff_2/lout')

wire n2081;
// (19, 22, 'lutff_7/lout')

wire n2082;
// (19, 13, 'lutff_6/lout')

wire n2083;
// (23, 11, 'lutff_1/lout')

wire n2084;
// (22, 17, 'lutff_1/lout')

wire n2085;
// (16, 16, 'lutff_7/lout')

wire n2086;
// (15, 13, 'lutff_5/lout')

wire n2087;
// (17, 13, 'lutff_0/lout')

wire n2088;
// (14, 16, 'lutff_4/out')

wire n2089;
// (16, 19, 'lutff_3/lout')

wire n2090;
// (13, 24, 'lutff_0/out')

wire n2091;
// (13, 24, 'lutff_0/lout')

wire n2092;
// (18, 17, 'lutff_5/out')

wire n2093;
// (20, 23, 'lutff_2/lout')

wire n2094;
// (10, 16, 'lutff_0/lout')

wire n2095;
// (13, 10, 'lutff_7/lout')

wire n2096;
// (18, 12, 'lutff_5/lout')

wire n2097;
// (14, 12, 'lutff_1/lout')

wire n2098;
// (19, 23, 'lutff_4/lout')

wire n2099;
// (19, 10, 'lutff_7/lout')

wire n2100;
// (22, 16, 'lutff_2/lout')

wire n2101;
// (26, 17, 'lutff_2/lout')

wire n2102;
// (14, 19, 'lutff_5/lout')

wire n2103;
// (17, 14, 'lutff_1/lout')

wire n2104;
// (19, 24, 'lutff_2/lout')

wire n2105;
// (11, 20, 'lutff_4/lout')

wire n2106;
// (16, 18, 'lutff_0/lout')

wire n2107;
// (15, 15, 'lutff_2/lout')

wire n2108;
// (20, 22, 'lutff_1/out')

wire n2109;
// (10, 19, 'lutff_1/lout')

wire n2110;
// (13, 22, 'lutff_7/lout')

wire n2111;
// (18, 15, 'lutff_4/out')

wire n2112;
// (14, 15, 'lutff_0/lout')

wire n2113;
// (19, 11, 'lutff_4/lout')

wire n2114;
// (22, 19, 'lutff_3/lout')

wire n2115;
// (17, 15, 'lutff_6/lout')

wire n2116;
// (11, 21, 'lutff_3/lout')

wire n2117;
// (16, 17, 'lutff_1/lout')

wire n2118;
// (22, 13, 'lutff_3/out')

wire n2119;
// (6, 8, 'lutff_1/lout')

wire n2120;
// (20, 21, 'lutff_0/lout')

wire n2121;
// (23, 13, 'lutff_4/lout')

wire n2122;
// (24, 14, 'lutff_4/lout')

wire n2123;
// (13, 12, 'lutff_1/lout')

wire n2124;
// (14, 21, 'lutff_6/lout')

wire n2125;
// (12, 20, 'lutff_0/lout')

wire n2126;
// (17, 11, 'lutff_3/out')

wire n2127;
// (19, 21, 'lutff_2/lout')

wire n2128;
// (23, 14, 'lutff_6/lout')

wire n2129;
// (24, 17, 'lutff_2/lout')

wire n2130;
// (21, 10, 'lutff_3/lout')

wire n2131;
// (12, 10, 'lutff_1/out')

wire n2132;
// (11, 18, 'lutff_2/lout')

wire n2133;
// (22, 12, 'lutff_0/lout')

wire n2134;
// (13, 16, 'lutff_4/lout')

wire n2135;
// (18, 18, 'lutff_0/lout')

wire n2136;
// (6, 11, 'lutff_0/lout')

// Carry-In for (6 11)
assign n112 = 1;

wire n2137;
// (23, 18, 'lutff_0/lout')

wire n2138;
// (14, 10, 'lutff_4/lout')

wire n2139;
// (16, 14, 'lutff_3/lout')

wire n2140;
// (5, 17, 'lutff_1/lout')

wire n2141;
// (13, 13, 'lutff_2/lout')

wire n2142;
// (14, 20, 'lutff_5/lout')

wire n2143;
// (17, 20, 'lutff_2/lout')

wire n2144;
// (19, 18, 'lutff_3/out')

wire n2145;
// (23, 15, 'lutff_5/lout')

wire n2146;
// (21, 16, 'lutff_5/out')

wire n2147;
// (21, 11, 'lutff_4/lout')

wire n2148;
// (18, 22, 'lutff_5/lout')

wire n2149;
// (17, 9, 'lutff_4/lout')

wire n2150;
// (11, 19, 'lutff_1/lout')

wire n2151;
// (10, 9, 'lutff_1/lout')

wire n2152;
// (22, 15, 'lutff_1/lout')

wire n2153;
// (13, 17, 'lutff_7/lout')

wire n2154;
// (18, 21, 'lutff_1/lout')

wire n2155;
// (19, 14, 'lutff_6/lout')

wire n2156;
// (16, 13, 'lutff_2/lout')

wire n2157;
// (5, 18, 'lutff_0/lout')

wire n2158;
// (10, 20, 'lutff_4/lout')

wire n2159;
// (18, 7, 'lutff_0/lout')

wire n2160;
// (21, 15, 'lutff_1/out')

wire n2161;
// (20, 25, 'lutff_1/lout')

wire n2162;
// (19, 19, 'lutff_0/lout')

wire n2163;
// (23, 12, 'lutff_4/lout')

wire n2164;
// (21, 17, 'lutff_6/lout')

wire n2165;
// (21, 12, 'lutff_5/lout')

wire n2166;
// (18, 25, 'lutff_4/lout')

wire n2167;
// (17, 10, 'lutff_5/lout')

wire n2168;
// (11, 16, 'lutff_0/out')

wire n2169;
// (22, 14, 'lutff_6/lout')

wire n2170;
// (13, 18, 'lutff_6/lout')

wire n2171;
// (18, 20, 'lutff_2/lout')

wire n2172;
// (23, 16, 'lutff_2/lout')

wire n2173;
// (11, 14, 'lutff_3/lout')

wire n2174;
// (16, 7, 'lutff_4/lout')

wire n2175;
// (19, 15, 'lutff_5/lout')

wire n2176;
// (16, 12, 'lutff_5/lout')

wire n2177;
// (15, 26, 'lutff_2/lout')

wire n2178;
// (12, 12, 'lutff_4/lout')

wire n2179;
// (14, 22, 'lutff_3/lout')

wire n2180;
// (17, 22, 'lutff_0/lout')

wire n2181;
// (17, 22, 'carry_in_mux')

// Carry-In for (17 22)
assign n2181 = 0;

wire n2182;
// (19, 16, 'lutff_1/lout')

wire n2183;
// (22, 10, 'lutff_3/lout')

wire n2184;
// (7, 11, 'lutff_6/lout')

wire n2185;
// (21, 18, 'lutff_7/lout')

wire n2186;
// (21, 13, 'lutff_6/lout')

wire n2187;
// (12, 15, 'lutff_6/lout')

wire n2188;
// (18, 24, 'lutff_7/lout')

wire n2189;
// (13, 19, 'lutff_1/lout')

wire n2190;
// (15, 21, 'lutff_0/lout')

wire n2191;
// (18, 23, 'lutff_3/lout')

wire n2192;
// (23, 17, 'lutff_5/lout')

wire n2193;
// (11, 15, 'lutff_0/lout')

wire n2194;
// (19, 12, 'lutff_4/lout')

wire n2195;
// (9, 19, 'lutff_2/lout')

wire n2196;
// (12, 19, 'lutff_5/lout')

wire n2197;
// (14, 17, 'lutff_2/lout')

wire n2198;
// (17, 12, 'lutff_6/lout')

wire n2199;
// (17, 23, 'lutff_7/lout')

wire n2200;
// (22, 21, 'lutff_1/lout')

wire n2201;
// (21, 19, 'lutff_0/out')

wire n2202;
// (13, 23, 'lutff_6/out')

wire n2203;
// (13, 23, 'lutff_6/lout')

wire n2204;
// (21, 14, 'lutff_7/lout')

wire n2205;
// (9, 16, 'lutff_4/lout')

wire n2206;
// (12, 14, 'lutff_5/lout')

wire n2207;
// (10, 10, 'lutff_4/lout')

wire n2208;
// (16, 23, 'lutff_3/lout')

wire n2209;
// (10, 17, 'lutff_6/out')

wire n2210;
// (10, 17, 'lutff_6/lout')

wire n2211;
// (13, 20, 'lutff_0/lout')

wire n2212;
// (15, 10, 'lutff_1/lout')

wire n2213;
// (20, 19, 'lutff_2/lout')

wire n2214;
// (11, 12, 'lutff_1/lout')

wire n2215;
// (17, 19, 'lutff_4/out')

wire n2216;
// (17, 19, 'lutff_4/lout')

wire n2217;
// (19, 13, 'lutff_3/lout')

wire n2218;
// (16, 10, 'lutff_7/lout')

wire n2219;
// (15, 24, 'lutff_0/lout')

// Carry-In for (15 24)
assign n1026 = 1;

wire n2220;
// (12, 18, 'lutff_6/lout')

wire n2221;
// (17, 13, 'lutff_5/lout')

wire n2222;
// (14, 16, 'lutff_1/lout')

wire n2223;
// (17, 16, 'lutff_6/lout')

wire n2224;
// (22, 20, 'lutff_2/out')

wire n2225;
// (10, 14, 'lutff_1/lout')

wire n2226;
// (21, 20, 'lutff_1/lout')

wire n2227;
// (13, 24, 'lutff_7/out')

wire n2228;
// (13, 24, 'lutff_7/lout')

wire n2229;
// (9, 17, 'lutff_7/lout')

wire n2230;
// (12, 13, 'lutff_4/lout')

wire n2231;
// (20, 12, 'lutff_0/lout')

wire n2232;
// (10, 13, 'lutff_5/lout')

wire n2233;
// (16, 22, 'lutff_0/lout')

wire n2234;
// (10, 16, 'lutff_5/lout')

wire n2235;
// (13, 21, 'lutff_3/lout')

wire n2236;
// (20, 18, 'lutff_1/lout')

wire n2237;
// (11, 13, 'lutff_6/lout')

wire n2238;
// (19, 10, 'lutff_2/lout')

wire n2239;
// (15, 25, 'lutff_7/lout')

wire n2240;
// (7, 13, 'lutff_5/lout')

wire n2241;
// (12, 17, 'lutff_7/lout')

wire n2242;
// (14, 19, 'lutff_0/lout')

wire n2243;
// (17, 14, 'lutff_4/lout')

wire n2244;
// (17, 17, 'lutff_5/out')

wire n2245;
// (22, 23, 'lutff_3/lout')

wire n2246;
// (21, 21, 'lutff_2/lout')

wire n2247;
// (16, 21, 'lutff_1/lout')

wire n2248;
// (10, 19, 'lutff_4/lout')

wire n2249;
// (13, 22, 'lutff_2/lout')

wire n2250;
// (6, 12, 'lutff_1/lout')

wire n2251;
// (20, 17, 'lutff_0/lout')

wire n2252;
// (23, 20, 'lutff_6/lout')

wire n2253;
// (11, 10, 'lutff_7/lout')

wire n2254;
// (19, 11, 'lutff_1/lout')

wire n2255;
// (12, 16, 'lutff_0/lout')

wire n2256;
// (17, 15, 'lutff_3/out')

wire n2257;
// (19, 25, 'lutff_2/lout')

wire n2258;
// (17, 18, 'lutff_4/out')

wire n2259;
// (17, 18, 'lutff_4/lout')

wire n2260;
// (22, 13, 'lutff_6/out')

wire n2261;
// (7, 15, 'lutff_2/lout')

wire n2262;
// (21, 22, 'lutff_3/lout')

wire n2263;
// (11, 22, 'lutff_2/lout')

wire n2264;
// (16, 15, 'lutff_7/lout')

wire n2265;
// (10, 15, 'lutff_7/lout')

wire n2266;
// (16, 20, 'lutff_6/lout')

wire n2267;
// (15, 18, 'lutff_5/lout')

wire n2268;
// (18, 14, 'lutff_0/out')

wire n2269;
// (20, 16, 'lutff_7/lout')

wire n2270;
// (12, 20, 'lutff_5/lout')

wire n2271;
// (11, 11, 'lutff_4/lout')

wire n2272;
// (22, 18, 'lutff_1/out')

wire n2273;
// (13, 9, 'lutff_2/lout')

wire n2274;
// (21, 10, 'lutff_6/lout')

wire n2275;
// (12, 23, 'lutff_1/out')

wire n2276;
// (12, 23, 'lutff_1/lout')

wire n2277;
// (17, 8, 'lutff_2/lout')

wire n2278;
// (19, 22, 'lutff_3/lout')

wire n2279;
// (22, 17, 'lutff_5/lout')

wire n2280;
// (16, 16, 'lutff_3/lout')

wire n2281;
// (22, 12, 'lutff_5/lout')

wire n2282;
// (20, 20, 'lutff_4/lout')

wire n2283;
// (16, 14, 'lutff_4/lout')

wire n2284;
// (16, 19, 'lutff_7/lout')

wire n2285;
// (15, 19, 'lutff_6/lout')

wire n2286;
// (15, 14, 'lutff_5/lout')

wire n2287;
// (18, 17, 'lutff_1/out')

wire n2288;
// (20, 23, 'lutff_6/lout')

wire n2289;
// (24, 16, 'lutff_2/lout')

wire n2290;
// (21, 11, 'lutff_1/lout')

wire n2291;
// (12, 22, 'lutff_2/out')

wire n2292;
// (12, 22, 'lutff_2/lout')

wire n2293;
// (19, 23, 'lutff_0/lout')

wire n2294;
// (22, 16, 'lutff_6/out')

wire n2295;
// (22, 15, 'lutff_4/lout')

wire n2296;
// (20, 11, 'lutff_5/lout')

wire n2297;
// (19, 24, 'lutff_6/lout')

wire n2298;
// (11, 20, 'lutff_0/lout')

wire n2299;
// (16, 13, 'lutff_5/lout')

wire n2300;
// (16, 18, 'lutff_4/lout')

wire n2301;
// (10, 20, 'lutff_1/lout')

wire n2302;
// (15, 16, 'lutff_7/lout')

wire n2303;
// (21, 15, 'lutff_6/lout')

wire n2304;
// (15, 15, 'lutff_6/lout')

wire n2305;
// (18, 16, 'lutff_2/lout')

wire n2306;
// (6, 9, 'lutff_6/lout')

wire n2307;
// (20, 22, 'lutff_5/lout')

wire n2308;
// (17, 24, 'lutff_1/out')

wire n2309;
// (17, 24, 'lutff_1/lout')

wire n2310;
// (24, 15, 'lutff_3/lout')

wire n2311;
// (21, 12, 'lutff_0/lout')

wire n2312;
// (12, 21, 'lutff_3/lout')

wire n2313;
// (17, 10, 'lutff_0/lout')

wire n2314;
// (19, 20, 'lutff_1/lout')

wire n2315;
// (22, 19, 'lutff_7/lout')

wire n2316;
// (22, 14, 'lutff_3/lout')

wire n2317;
// (23, 16, 'lutff_5/lout')

wire n2318;
// (11, 14, 'lutff_6/lout')

wire n2319;
// (16, 12, 'lutff_2/out')

wire n2320;
// (16, 17, 'lutff_5/lout')

wire n2321;
// (13, 15, 'lutff_1/lout')

wire n2322;
// (15, 17, 'lutff_0/lout')

wire n2323;
// (15, 12, 'lutff_7/lout')

wire n2324;
// (18, 19, 'lutff_3/lout')

wire n2325;
// (20, 21, 'lutff_4/lout')

wire n2326;
// (24, 14, 'lutff_0/lout')

wire n2327;
// (13, 12, 'lutff_5/lout')

wire n2328;
// (21, 13, 'lutff_3/lout')

wire n2329;
// (19, 21, 'lutff_6/lout')

wire n2330;
// (24, 17, 'lutff_6/lout')

wire n2331;
// (15, 21, 'lutff_5/lout')

wire n2332;
// (20, 9, 'lutff_7/lout')

wire n2333;
// (23, 17, 'lutff_2/lout')

wire n2334;
// (11, 15, 'lutff_5/lout')

wire n2335;
// (11, 18, 'lutff_6/lout')

wire n2336;
// (16, 11, 'lutff_3/lout')

wire n2337;
// (13, 16, 'lutff_0/lout')

wire n2338;
// (15, 22, 'lutff_1/out')

wire n2339;
// (15, 22, 'lutff_1/lout')

wire n2340;
// (18, 9, 'lutff_5/lout')

wire n2341;
// (18, 18, 'lutff_4/lout')

wire n2342;
// (6, 11, 'lutff_4/lout')

wire n2343;
// (14, 10, 'lutff_0/lout')

wire n2344;
// (19, 17, 'lutff_3/lout')

wire n2345;
// (22, 21, 'lutff_4/lout')

wire n2346;
// (24, 13, 'lutff_1/lout')

wire n2347;
// (13, 13, 'lutff_6/lout')

wire n2348;
// (21, 14, 'lutff_2/lout')

wire n2349;
// (9, 16, 'lutff_3/lout')

wire n2350;
// (14, 20, 'lutff_1/lout')

wire n2351;
// (19, 18, 'lutff_7/lout')

wire n2352;
// (10, 10, 'lutff_1/lout')

wire n2353;
// (16, 23, 'lutff_6/lout')

wire n2354;
// (21, 16, 'lutff_1/out')

wire n2355;
// (15, 10, 'lutff_4/lout')

wire n2356;
// (11, 12, 'lutff_4/lout')

wire n2357;
// (11, 19, 'lutff_5/lout')

wire n2358;
// (16, 10, 'lutff_0/lout')

wire n2359;
// (9, 12, 'lutff_5/lout')

wire n2360;
// (18, 21, 'lutff_5/lout')

wire n2361;
// (19, 14, 'lutff_2/lout')

wire n2362;
// (22, 20, 'lutff_7/lout')

wire n2363;
// (16, 24, 'lutff_4/lout')

wire n2364;
// (9, 17, 'lutff_0/lout')

wire n2365;
// (20, 12, 'lutff_5/lout')

wire n2366;
// (19, 19, 'lutff_4/lout')

wire n2367;
// (10, 13, 'lutff_0/lout')

// Carry-In for (10 13)
assign n305 = 1;

wire n2368;
// (16, 22, 'lutff_5/lout')

wire n2369;
// (22, 11, 'lutff_0/lout')

wire n2370;
// (21, 17, 'lutff_2/lout')

wire n2371;
// (20, 15, 'lutff_1/lout')

wire n2372;
// (11, 13, 'lutff_3/lout')

wire n2373;
// (11, 16, 'lutff_4/lout')

wire n2374;
// (16, 9, 'lutff_1/lout')

wire n2375;
// (13, 18, 'lutff_2/lout')

wire n2376;
// (15, 20, 'lutff_3/lout')

wire n2377;
// (18, 20, 'lutff_6/lout')

wire n2378;
// (16, 7, 'lutff_0/lout')

wire n2379;
// (16, 7, 'carry_in_mux')

// Carry-In for (16 7)
assign n2379 = 0;

wire n2380;
// (19, 15, 'lutff_1/out')

wire n2381;
// (22, 23, 'lutff_6/lout')

wire n2382;
// (24, 22, 'lutff_4/lout')

wire n2383;
// (9, 18, 'lutff_1/lout')

wire n2384;
// (12, 12, 'lutff_0/lout')

wire n2385;
// (19, 16, 'lutff_5/lout')

wire n2386;
// (16, 21, 'lutff_4/lout')

wire n2387;
// (16, 26, 'lutff_5/lout')

wire n2388;
// (21, 18, 'lutff_3/out')

wire n2389;
// (15, 7, 'lutff_7/lout')

wire n2390;
// (18, 24, 'lutff_3/out')

wire n2391;
// (20, 14, 'lutff_2/lout')

wire n2392;
// (23, 20, 'lutff_1/lout')

wire n2393;
// (11, 10, 'lutff_2/out')

wire n2394;
// (9, 14, 'lutff_7/lout')

wire n2395;
// (13, 19, 'lutff_5/lout')

wire n2396;
// (18, 23, 'lutff_7/lout')

wire n2397;
// (14, 18, 'lutff_4/lout')

wire n2398;
// (14, 7, 'lutff_3/lout')

wire n2399;
// (19, 12, 'lutff_0/lout')

wire n2400;
// (22, 22, 'lutff_1/lout')

wire n2401;
// (12, 19, 'lutff_1/lout')

wire n2402;
// (17, 12, 'lutff_2/lout')

wire n2403;
// (10, 15, 'lutff_2/lout')

wire n2404;
// (16, 20, 'lutff_3/lout')

wire n2405;
// (21, 19, 'lutff_4/out')

wire n2406;
// (13, 23, 'lutff_2/out')

wire n2407;
// (13, 23, 'lutff_2/lout')

wire n2408;
// (15, 9, 'lutff_1/lout')

wire n2409;
// (18, 14, 'lutff_5/lout')

wire n2410;
// (20, 13, 'lutff_3/out')

wire n2411;
// (11, 11, 'lutff_1/lout')

wire n2412;
// (22, 18, 'lutff_6/lout')

wire n2413;
// (10, 17, 'lutff_2/lout')

wire n2414;
// (9, 15, 'lutff_0/lout')

wire n2415;
// (13, 20, 'lutff_4/lout')

wire n2416;
// (18, 13, 'lutff_1/lout')

wire n2417;
// (14, 13, 'lutff_5/lout')

wire n2418;
// (19, 22, 'lutff_6/lout')

wire n2419;
// (17, 19, 'lutff_0/out')

wire n2420;
// (17, 19, 'lutff_0/lout')

wire n2421;
// (19, 13, 'lutff_7/lout')

wire n2422;
// (22, 17, 'lutff_0/out')

wire n2423;
// (15, 13, 'lutff_6/lout')

wire n2424;
// (12, 18, 'lutff_2/lout')

wire n2425;
// (14, 16, 'lutff_5/lout')

wire n2426;
// (17, 13, 'lutff_1/out')

wire n2427;
// (16, 19, 'lutff_2/lout')

wire n2428;
// (21, 20, 'lutff_5/lout')

wire n2429;
// (13, 24, 'lutff_3/out')

wire n2430;
// (13, 24, 'lutff_3/lout')

wire n2431;
// (18, 17, 'lutff_4/out')

wire n2432;
// (18, 26, 'lutff_5/lout')

wire n2433;
// (10, 16, 'lutff_1/lout')

wire n2434;
// (13, 21, 'lutff_7/lout')

wire n2435;
// (18, 12, 'lutff_2/lout')

wire n2436;
// (14, 12, 'lutff_6/lout')

wire n2437;
// (19, 23, 'lutff_5/lout')

wire n2438;
// (19, 10, 'lutff_6/lout')

wire n2439;
// (22, 16, 'lutff_3/out')

wire n2440;
// (12, 17, 'lutff_3/lout')

wire n2441;
// (14, 19, 'lutff_4/lout')

wire n2442;
// (17, 14, 'lutff_0/out')

wire n2443;
// (19, 24, 'lutff_1/lout')

wire n2444;
// (16, 18, 'lutff_1/lout')

wire n2445;
// (21, 21, 'lutff_6/lout')

wire n2446;
// (13, 25, 'lutff_0/lout')

wire n2447;
// (15, 15, 'lutff_3/lout')

wire n2448;
// (10, 19, 'lutff_0/lout')

wire n2449;
// (13, 11, 'lutff_1/lout')

wire n2450;
// (13, 22, 'lutff_6/lout')

wire n2451;
// (18, 15, 'lutff_3/lout')

wire n2452;
// (14, 15, 'lutff_7/lout')

wire n2453;
// (19, 20, 'lutff_4/lout')

wire n2454;
// (19, 11, 'lutff_5/lout')

wire n2455;
// (22, 19, 'lutff_2/lout')

wire n2456;
// (17, 15, 'lutff_7/lout')

wire n2457;
// (16, 17, 'lutff_0/lout')

wire n2458;
// (22, 13, 'lutff_2/lout')

wire n2459;
// (15, 12, 'lutff_2/lout')

wire n2460;
// (18, 19, 'lutff_6/lout')

wire n2461;
// (23, 13, 'lutff_5/lout')

wire n2462;
// (24, 14, 'lutff_5/lout')

wire n2463;
// (9, 10, 'lutff_3/lout')

wire n2464;
// (13, 12, 'lutff_0/out')

wire n2465;
// (13, 12, 'lutff_0/lout')

wire n2466;
// (13, 12, 'carry_in_mux')

// Carry-In for (13 12)
assign n2466 = 0;

wire n2467;
// (15, 18, 'lutff_1/lout')

wire n2468;
// (14, 14, 'lutff_0/lout')

wire n2469;
// (17, 11, 'lutff_4/lout')

wire n2470;
// (19, 21, 'lutff_3/lout')

wire n2471;
// (23, 14, 'lutff_1/lout')

wire n2472;
// (24, 17, 'lutff_1/lout')

wire n2473;
// (21, 10, 'lutff_2/lout')

wire n2474;
// (12, 23, 'lutff_5/out')

wire n2475;
// (12, 23, 'lutff_5/lout')

wire n2476;
// (22, 12, 'lutff_1/lout')

wire n2477;
// (13, 16, 'lutff_7/lout')

wire n2478;
// (7, 12, 'lutff_7/lout')

wire n2479;
// (18, 18, 'lutff_1/out')

wire n2480;
// (20, 20, 'lutff_0/lout')

wire n2481;
// (23, 18, 'lutff_3/lout')

wire n2482;
// (14, 10, 'lutff_5/lout')

wire n2483;
// (16, 14, 'lutff_0/lout')

wire n2484;
// (5, 17, 'lutff_6/lout')

wire n2485;
// (13, 13, 'lutff_3/lout')

wire n2486;
// (17, 20, 'lutff_5/lout')

wire n2487;
// (19, 18, 'lutff_2/lout')

wire n2488;
// (23, 15, 'lutff_2/lout')

wire n2489;
// (21, 16, 'lutff_4/lout')

wire n2490;
// (21, 11, 'lutff_5/lout')

wire n2491;
// (18, 22, 'lutff_6/lout')

wire n2492;
// (12, 22, 'lutff_6/out')

wire n2493;
// (12, 22, 'lutff_6/lout')

wire n2494;
// (10, 9, 'lutff_0/lout')

wire n2495;
// (22, 15, 'lutff_0/lout')

wire n2496;
// (13, 17, 'lutff_4/lout')

wire n2497;
// (18, 21, 'lutff_0/lout')

wire n2498;
// (20, 11, 'lutff_1/lout')

wire n2499;
// (16, 13, 'lutff_1/lout')

wire n2500;
// (5, 18, 'lutff_7/lout')

wire n2501;
// (10, 20, 'lutff_5/lout')

wire n2502;
// (15, 16, 'lutff_3/lout')

wire n2503;
// (21, 15, 'lutff_2/lout')

wire n2504;
// (20, 25, 'lutff_0/lout')

wire n2505;
// (17, 21, 'lutff_6/lout')

wire n2506;
// (19, 19, 'lutff_1/lout')

wire n2507;
// (17, 24, 'lutff_5/out')

wire n2508;
// (17, 24, 'lutff_5/lout')

wire n2509;
// (23, 12, 'lutff_3/lout')

wire n2510;
// (21, 17, 'lutff_7/lout')

wire n2511;
// (21, 12, 'lutff_4/lout')

wire n2512;
// (12, 21, 'lutff_7/lout')

wire n2513;
// (17, 10, 'lutff_4/lout')

wire n2514;
// (22, 14, 'lutff_7/lout')

wire n2515;
// (13, 18, 'lutff_5/lout')

wire n2516;
// (23, 16, 'lutff_1/lout')

wire n2517;
// (11, 14, 'lutff_2/lout')

wire n2518;
// (5, 19, 'lutff_0/lout')

wire n2519;
// (22, 24, 'lutff_0/lout')

wire n2520;
// (15, 17, 'lutff_4/lout')

wire n2521;
// (20, 24, 'lutff_7/lout')

wire n2522;
// (17, 22, 'lutff_7/lout')

wire n2523;
// (14, 11, 'lutff_3/lout')

wire n2524;
// (19, 16, 'lutff_0/lout')

wire n2525;
// (22, 10, 'lutff_4/lout')

wire n2526;
// (21, 18, 'lutff_6/out')

wire n2527;
// (21, 13, 'lutff_7/lout')

wire n2528;
// (12, 15, 'lutff_1/lout')

wire n2529;
// (15, 7, 'lutff_0/lout')

wire n2530;
// (18, 24, 'lutff_4/out')

wire n2531;
// (13, 19, 'lutff_2/lout')

wire n2532;
// (15, 21, 'lutff_1/lout')

wire n2533;
// (18, 23, 'lutff_2/lout')

wire n2534;
// (23, 17, 'lutff_6/out')

wire n2535;
// (11, 15, 'lutff_1/lout')

wire n2536;
// (16, 11, 'lutff_7/lout')

wire n2537;
// (5, 20, 'lutff_1/lout')

wire n2538;
// (15, 22, 'lutff_5/out')

wire n2539;
// (15, 22, 'lutff_5/lout')

wire n2540;
// (18, 9, 'lutff_1/lout')

wire n2541;
// (12, 19, 'lutff_4/lout')

wire n2542;
// (17, 23, 'lutff_0/lout')

wire n2543;
// (22, 21, 'lutff_0/lout')

wire n2544;
// (21, 19, 'lutff_1/out')

wire n2545;
// (13, 23, 'lutff_7/out')

wire n2546;
// (13, 23, 'lutff_7/lout')

wire n2547;
// (21, 14, 'lutff_6/out')

wire n2548;
// (9, 16, 'lutff_7/lout')

wire n2549;
// (12, 14, 'lutff_2/lout')

wire n2550;
// (10, 10, 'lutff_5/out')

wire n2551;
// (10, 10, 'lutff_5/lout')

wire n2552;
// (16, 23, 'lutff_2/lout')

wire n2553;
// (13, 20, 'lutff_3/lout')

wire n2554;
// (15, 10, 'lutff_0/lout')

wire n2555;
// (20, 19, 'lutff_5/lout')

wire n2556;
// (11, 12, 'lutff_0/lout')

wire n2557;
// (17, 19, 'lutff_5/out')

wire n2558;
// (17, 19, 'lutff_5/lout')

wire n2559;
// (16, 10, 'lutff_4/lout')

wire n2560;
// (9, 12, 'lutff_1/lout')

wire n2561;
// (15, 24, 'lutff_7/lout')

wire n2562;
// (12, 18, 'lutff_7/lout')

wire n2563;
// (17, 16, 'lutff_1/lout')

wire n2564;
// (22, 20, 'lutff_3/out')

wire n2565;
// (10, 14, 'lutff_2/lout')

wire n2566;
// (16, 24, 'lutff_0/lout')

wire n2567;
// (21, 20, 'lutff_0/lout')

wire n2568;
// (13, 24, 'lutff_6/out')

wire n2569;
// (13, 24, 'lutff_6/lout')

wire n2570;
// (12, 13, 'lutff_3/lout')

wire n2571;
// (20, 12, 'lutff_1/lout')

wire n2572;
// (10, 13, 'lutff_4/lout')

wire n2573;
// (16, 22, 'lutff_1/lout')

wire n2574;
// (13, 21, 'lutff_0/lout')

wire n2575;
// (20, 18, 'lutff_6/lout')

wire n2576;
// (20, 15, 'lutff_5/lout')

wire n2577;
// (11, 13, 'lutff_7/lout')

wire n2578;
// (13, 7, 'lutff_1/out')

wire n2579;
// (15, 25, 'lutff_0/lout')

wire n2580;
// (15, 20, 'lutff_7/lout')

wire n2581;
// (18, 11, 'lutff_3/lout')

wire n2582;
// (12, 17, 'lutff_6/lout')

wire n2583;
// (17, 17, 'lutff_2/lout')

wire n2584;
// (22, 23, 'lutff_2/lout')

wire n2585;
// (11, 9, 'lutff_4/lout')

wire n2586;
// (16, 21, 'lutff_0/lout')

wire n2587;
// (13, 22, 'lutff_1/lout')

wire n2588;
// (20, 17, 'lutff_7/lout')

wire n2589;
// (20, 14, 'lutff_6/lout')

wire n2590;
// (23, 20, 'lutff_5/lout')

wire n2591;
// (14, 18, 'lutff_0/lout')

// Carry-In for (14 18)
assign n827 = 1;

wire n2592;
// (17, 18, 'lutff_3/out')

wire n2593;
// (17, 18, 'lutff_3/lout')

wire n2594;
// (21, 22, 'lutff_2/lout')

wire n2595;
// (11, 22, 'lutff_5/lout')

wire n2596;
// (10, 15, 'lutff_6/lout')

wire n2597;
// (16, 20, 'lutff_7/lout')

wire n2598;
// (21, 24, 'lutff_1/lout')

wire n2599;
// (15, 18, 'lutff_4/lout')

wire n2600;
// (18, 14, 'lutff_1/lout')

wire n2601;
// (20, 16, 'lutff_0/lout')

wire n2602;
// (12, 20, 'lutff_6/lout')

wire n2603;
// (20, 13, 'lutff_7/lout')

wire n2604;
// (11, 11, 'lutff_5/lout')

wire n2605;
// (22, 18, 'lutff_2/lout')

wire n2606;
// (9, 15, 'lutff_4/lout')

wire n2607;
// (12, 23, 'lutff_0/out')

wire n2608;
// (12, 23, 'lutff_0/lout')

wire n2609;
// (14, 13, 'lutff_1/lout')

wire n2610;
// (19, 22, 'lutff_2/lout')

wire n2611;
// (22, 17, 'lutff_4/out')

wire n2612;
// (16, 16, 'lutff_4/lout')

wire n2613;
// (7, 12, 'lutff_2/lout')

wire n2614;
// (15, 13, 'lutff_2/lout')

wire n2615;
// (20, 20, 'lutff_5/lout')

wire n2616;
// (16, 19, 'lutff_6/lout')

wire n2617;
// (15, 19, 'lutff_7/lout')

wire n2618;
// (18, 17, 'lutff_0/lout')

wire n2619;
// (15, 14, 'lutff_4/lout')

wire n2620;
// (19, 9, 'lutff_0/lout')

wire n2621;
// (21, 11, 'lutff_2/lout')

wire n2622;
// (18, 12, 'lutff_6/lout')

wire n2623;
// (12, 22, 'lutff_3/out')

wire n2624;
// (12, 22, 'lutff_3/lout')

wire n2625;
// (14, 12, 'lutff_2/lout')

wire n2626;
// (19, 23, 'lutff_1/lout')

wire n2627;
// (22, 16, 'lutff_7/lout')

wire n2628;
// (20, 11, 'lutff_4/lout')

wire n2629;
// (19, 24, 'lutff_5/lout')

wire n2630;
// (11, 20, 'lutff_7/lout')

wire n2631;
// (16, 13, 'lutff_4/lout')

wire n2632;
// (16, 18, 'lutff_5/lout')

wire n2633;
// (21, 15, 'lutff_7/lout')

wire n2634;
// (15, 15, 'lutff_7/lout')

wire n2635;
// (18, 16, 'lutff_3/lout')

wire n2636;
// (20, 22, 'lutff_2/lout')

wire n2637;
// (17, 24, 'lutff_0/out')

wire n2638;
// (17, 24, 'lutff_0/lout')

wire n2639;
// (24, 15, 'lutff_2/lout')

wire n2640;
// (13, 11, 'lutff_5/lout')

wire n2641;
// (21, 12, 'lutff_3/lout')

wire n2642;
// (12, 21, 'lutff_2/lout')

wire n2643;
// (19, 20, 'lutff_0/lout')

wire n2644;
// (22, 19, 'lutff_6/lout')

wire n2645;
// (23, 16, 'lutff_4/lout')

wire n2646;
// (11, 21, 'lutff_0/lout')

wire n2647;
// (16, 12, 'lutff_3/out')

wire n2648;
// (16, 17, 'lutff_4/lout')

wire n2649;
// (13, 15, 'lutff_2/lout')

wire n2650;
// (15, 17, 'lutff_1/lout')

wire n2651;
// (18, 19, 'lutff_2/lout')

wire n2652;
// (20, 21, 'lutff_3/lout')

wire n2653;
// (17, 25, 'lutff_3/lout')

wire n2654;
// (23, 13, 'lutff_1/lout')

wire n2655;
// (24, 14, 'lutff_1/lout')

wire n2656;
// (13, 12, 'lutff_4/lout')

wire n2657;
// (21, 13, 'lutff_0/lout')

wire n2658;
// (17, 11, 'lutff_0/lout')

wire n2659;
// (19, 21, 'lutff_7/lout')

wire n2660;
// (11, 17, 'lutff_5/lout')

wire n2661;
// (23, 14, 'lutff_5/lout')

wire n2662;
// (24, 17, 'lutff_5/lout')

wire n2663;
// (15, 21, 'lutff_6/lout')

wire n2664;
// (12, 10, 'lutff_2/out')

wire n2665;
// (23, 17, 'lutff_3/out')

wire n2666;
// (11, 18, 'lutff_1/lout')

wire n2667;
// (16, 11, 'lutff_2/lout')

wire n2668;
// (13, 16, 'lutff_3/lout')

wire n2669;
// (15, 22, 'lutff_0/out')

wire n2670;
// (15, 22, 'lutff_0/lout')

wire n2671;
// (18, 9, 'lutff_4/lout')

wire n2672;
// (18, 18, 'lutff_5/out')

wire n2673;
// (6, 11, 'lutff_3/lout')

wire n2674;
// (14, 10, 'lutff_1/lout')

wire n2675;
// (19, 17, 'lutff_4/out')

wire n2676;
// (22, 21, 'lutff_7/lout')

wire n2677;
// (5, 17, 'lutff_2/lout')

wire n2678;
// (24, 13, 'lutff_0/lout')

wire n2679;
// (21, 14, 'lutff_1/lout')

wire n2680;
// (9, 16, 'lutff_2/lout')

wire n2681;
// (14, 20, 'lutff_6/lout')

wire n2682;
// (14, 9, 'lutff_5/lout')

wire n2683;
// (17, 20, 'lutff_1/lout')

wire n2684;
// (19, 18, 'lutff_6/lout')

wire n2685;
// (10, 10, 'lutff_2/lout')

wire n2686;
// (23, 15, 'lutff_6/lout')

wire n2687;
// (21, 16, 'lutff_0/lout')

wire n2688;
// (15, 10, 'lutff_7/lout')

wire n2689;
// (12, 9, 'lutff_3/lout')

wire n2690;
// (11, 19, 'lutff_2/lout')

wire n2691;
// (9, 12, 'lutff_4/lout')

wire n2692;
// (13, 17, 'lutff_0/lout')

wire n2693;
// (18, 21, 'lutff_4/lout')

wire n2694;
// (19, 14, 'lutff_5/lout')

wire n2695;
// (22, 20, 'lutff_4/lout')

wire n2696;
// (10, 14, 'lutff_7/lout')

wire n2697;
// (5, 18, 'lutff_3/lout')

wire n2698;
// (16, 24, 'lutff_5/lout')

wire n2699;
// (9, 17, 'lutff_1/lout')

wire n2700;
// (14, 23, 'lutff_7/lout')

wire n2701;
// (20, 12, 'lutff_6/lout')

wire n2702;
// (19, 19, 'lutff_5/lout')

wire n2703;
// (10, 13, 'lutff_3/lout')

wire n2704;
// (23, 12, 'lutff_7/lout')

wire n2705;
// (21, 17, 'lutff_3/lout')

wire n2706;
// (15, 11, 'lutff_4/lout')

wire n2707;
// (18, 25, 'lutff_3/lout')

wire n2708;
// (20, 15, 'lutff_0/lout')

wire n2709;
// (11, 16, 'lutff_3/lout')

wire n2710;
// (16, 9, 'lutff_0/lout')

wire n2711;
// (13, 18, 'lutff_1/lout')

wire n2712;
// (15, 20, 'lutff_2/lout')

wire n2713;
// (18, 20, 'lutff_7/lout')

wire n2714;
// (16, 7, 'lutff_3/lout')

wire n2715;
// (19, 15, 'lutff_6/out')

wire n2716;
// (22, 23, 'lutff_5/lout')

wire n2717;
// (15, 26, 'lutff_1/lout')

wire n2718;
// (9, 18, 'lutff_0/lout')

wire n2719;
// (12, 12, 'lutff_1/lout')

wire n2720;
// (14, 22, 'lutff_0/lout')

wire n2721;
// (17, 22, 'lutff_3/lout')

wire n2722;
// (14, 11, 'lutff_7/lout')

wire n2723;
// (19, 16, 'lutff_4/lout')

wire n2724;
// (22, 10, 'lutff_0/out')

wire n2725;
// (22, 10, 'lutff_0/lout')

wire n2726;
// (22, 10, 'carry_in_mux')

// Carry-In for (22 10)
assign n2726 = 0;

wire n2727;
// (21, 18, 'lutff_2/lout')

wire n2728;
// (12, 15, 'lutff_5/lout')

wire n2729;
// (15, 7, 'lutff_4/lout')

wire n2730;
// (20, 14, 'lutff_3/out')

wire n2731;
// (23, 20, 'lutff_0/lout')

wire n2732;
// (13, 19, 'lutff_6/lout')

wire n2733;
// (18, 23, 'lutff_6/lout')

wire n2734;
// (14, 18, 'lutff_5/lout')

wire n2735;
// (14, 7, 'lutff_2/lout')

wire n2736;
// (19, 12, 'lutff_7/lout')

wire n2737;
// (12, 19, 'lutff_0/lout')

wire n2738;
// (14, 17, 'lutff_1/lout')

wire n2739;
// (17, 12, 'lutff_5/lout')

wire n2740;
// (17, 23, 'lutff_4/lout')

wire n2741;
// (10, 15, 'lutff_1/lout')

wire n2742;
// (21, 19, 'lutff_5/out')

wire n2743;
// (13, 23, 'lutff_3/out')

wire n2744;
// (13, 23, 'lutff_3/lout')

wire n2745;
// (18, 14, 'lutff_6/lout')

wire n2746;
// (15, 9, 'lutff_2/lout')

wire n2747;
// (12, 14, 'lutff_6/lout')

wire n2748;
// (20, 13, 'lutff_2/lout')

wire n2749;
// (10, 17, 'lutff_5/lout')

wire n2750;
// (9, 15, 'lutff_1/lout')

wire n2751;
// (13, 20, 'lutff_7/lout')

wire n2752;
// (18, 13, 'lutff_0/out')

wire n2753;
// (20, 19, 'lutff_1/lout')

wire n2754;
// (14, 13, 'lutff_4/lout')

wire n2755;
// (17, 19, 'lutff_1/out')

wire n2756;
// (17, 19, 'lutff_1/lout')

wire n2757;
// (19, 13, 'lutff_0/lout')

wire n2758;
// (22, 17, 'lutff_3/lout')

wire n2759;
// (15, 24, 'lutff_3/lout')

wire n2760;
// (21, 23, 'lutff_2/lout')

wire n2761;
// (15, 13, 'lutff_7/lout')

wire n2762;
// (12, 18, 'lutff_3/lout')

wire n2763;
// (14, 16, 'lutff_2/lout')

wire n2764;
// (17, 13, 'lutff_6/out')

wire n2765;
// (17, 16, 'lutff_5/out')

wire n2766;
// (21, 20, 'lutff_4/lout')

wire n2767;
// (13, 24, 'lutff_2/out')

wire n2768;
// (13, 24, 'lutff_2/lout')

wire n2769;
// (15, 14, 'lutff_3/lout')

wire n2770;
// (18, 17, 'lutff_7/lout')

wire n2771;
// (12, 13, 'lutff_7/lout')

wire n2772;
// (10, 16, 'lutff_6/lout')

wire n2773;
// (18, 12, 'lutff_3/lout')

wire n2774;
// (20, 18, 'lutff_2/lout')

wire n2775;
// (19, 10, 'lutff_1/lout')

wire n2776;
// (22, 16, 'lutff_0/lout')

wire n2777;
// (15, 25, 'lutff_4/lout')

wire n2778;
// (12, 17, 'lutff_2/lout')

wire n2779;
// (14, 19, 'lutff_3/lout')

wire n2780;
// (17, 14, 'lutff_7/lout')

wire n2781;
// (19, 24, 'lutff_0/lout')

// Carry-In for (19 24)
assign n1525 = 1;

wire n2782;
// (17, 17, 'lutff_6/lout')

wire n2783;
// (21, 21, 'lutff_7/lout')

wire n2784;
// (15, 15, 'lutff_0/lout')

wire n2785;
// (18, 16, 'lutff_4/lout')

wire n2786;
// (10, 19, 'lutff_7/lout')

wire n2787;
// (13, 11, 'lutff_2/lout')

wire n2788;
// (13, 22, 'lutff_5/lout')

wire n2789;
// (18, 15, 'lutff_2/out')

wire n2790;
// (6, 12, 'lutff_2/lout')

wire n2791;
// (20, 17, 'lutff_3/lout')

wire n2792;
// (14, 15, 'lutff_6/lout')

wire n2793;
// (19, 11, 'lutff_2/lout')

wire n2794;
// (22, 19, 'lutff_1/lout')

wire n2795;
// (12, 16, 'lutff_5/lout')

wire n2796;
// (17, 15, 'lutff_0/out')

wire n2797;
// (17, 18, 'lutff_7/out')

wire n2798;
// (17, 18, 'lutff_7/lout')

wire n2799;
// (22, 13, 'lutff_5/lout')

wire n2800;
// (15, 12, 'lutff_1/lout')

wire n2801;
// (18, 19, 'lutff_5/lout')

wire n2802;
// (11, 22, 'lutff_1/lout')

wire n2803;
// (16, 15, 'lutff_2/lout')

wire n2804;
// (10, 18, 'lutff_0/lout')

wire n2805;
// (13, 12, 'lutff_3/lout')

wire n2806;
// (15, 18, 'lutff_0/lout')

wire n2807;
// (20, 16, 'lutff_4/lout')

wire n2808;
// (12, 20, 'lutff_2/lout')

wire n2809;
// (14, 14, 'lutff_1/lout')

wire n2810;
// (17, 11, 'lutff_5/lout')

wire n2811;
// (19, 8, 'lutff_3/lout')

wire n2812;
// (23, 14, 'lutff_0/lout')

wire n2813;
// (24, 17, 'lutff_0/lout')

wire n2814;
// (21, 10, 'lutff_1/lout')

wire n2815;
// (12, 10, 'lutff_7/lout')

wire n2816;
// (12, 23, 'lutff_4/out')

wire n2817;
// (12, 23, 'lutff_4/lout')

wire n2818;
// (17, 8, 'lutff_1/lout')

wire n2819;
// (16, 16, 'lutff_0/lout')

wire n2820;
// (22, 12, 'lutff_6/lout')

wire n2821;
// (13, 16, 'lutff_6/lout')

wire n2822;
// (18, 18, 'lutff_2/lout')

wire n2823;
// (20, 20, 'lutff_1/lout')

wire n2824;
// (23, 18, 'lutff_2/lout')

wire n2825;
// (16, 14, 'lutff_1/lout')

wire n2826;
// (5, 17, 'lutff_7/lout')

wire n2827;
// (13, 13, 'lutff_0/lout')

wire n2828;
// (15, 19, 'lutff_3/lout')

wire n2829;
// (20, 23, 'lutff_5/lout')

wire n2830;
// (14, 9, 'lutff_0/lout')

wire n2831;
// (17, 20, 'lutff_4/lout')

wire n2832;
// (23, 15, 'lutff_3/lout')

wire n2833;
// (21, 16, 'lutff_7/lout')

wire n2834;
// (21, 11, 'lutff_6/lout')

wire n2835;
// (18, 22, 'lutff_7/lout')

wire n2836;
// (12, 22, 'lutff_7/out')

wire n2837;
// (12, 22, 'lutff_7/lout')

wire n2838;
// (10, 9, 'lutff_3/lout')

wire n2839;
// (22, 15, 'lutff_7/lout')

wire n2840;
// (13, 17, 'lutff_5/lout')

wire n2841;
// (18, 21, 'lutff_3/lout')

wire n2842;
// (20, 11, 'lutff_0/lout')

wire n2843;
// (23, 19, 'lutff_1/lout')

wire n2844;
// (11, 20, 'lutff_3/lout')

wire n2845;
// (16, 13, 'lutff_0/lout')

wire n2846;
// (5, 18, 'lutff_6/lout')

wire n2847;
// (10, 20, 'lutff_2/lout')

wire n2848;
// (15, 16, 'lutff_2/lout')

wire n2849;
// (21, 15, 'lutff_3/out')

wire n2850;
// (20, 25, 'lutff_7/lout')

wire n2851;
// (20, 22, 'lutff_6/lout')

wire n2852;
// (17, 24, 'lutff_4/out')

wire n2853;
// (17, 24, 'lutff_4/lout')

wire n2854;
// (23, 12, 'lutff_2/lout')

wire n2855;
// (7, 10, 'lutff_7/lout')

wire n2856;
// (21, 17, 'lutff_4/lout')

wire n2857;
// (21, 12, 'lutff_7/lout')

wire n2858;
// (18, 25, 'lutff_6/lout')

wire n2859;
// (12, 21, 'lutff_6/lout')

wire n2860;
// (22, 14, 'lutff_0/lout')

wire n2861;
// (13, 18, 'lutff_4/lout')

wire n2862;
// (18, 20, 'lutff_0/out')

wire n2863;
// (20, 10, 'lutff_3/lout')

wire n2864;
// (23, 16, 'lutff_0/lout')

wire n2865;
// (11, 14, 'lutff_5/lout')

wire n2866;
// (16, 12, 'lutff_7/lout')

wire n2867;
// (5, 19, 'lutff_1/lout')

wire n2868;
// (22, 24, 'lutff_1/lout')

wire n2869;
// (15, 17, 'lutff_5/lout')

wire n2870;
// (12, 12, 'lutff_6/lout')

wire n2871;
// (20, 21, 'lutff_7/lout')

wire n2872;
// (17, 22, 'lutff_6/lout')

wire n2873;
// (14, 11, 'lutff_2/lout')

wire n2874;
// (22, 10, 'lutff_5/lout')

wire n2875;
// (21, 18, 'lutff_5/lout')

wire n2876;
// (21, 13, 'lutff_4/lout')

wire n2877;
// (12, 15, 'lutff_0/lout')

wire n2878;
// (18, 24, 'lutff_5/lout')

wire n2879;
// (11, 17, 'lutff_1/lout')

wire n2880;
// (13, 19, 'lutff_3/lout')

wire n2881;
// (15, 21, 'lutff_2/lout')

wire n2882;
// (18, 23, 'lutff_1/lout')

wire n2883;
// (23, 17, 'lutff_7/lout')

wire n2884;
// (11, 15, 'lutff_6/lout')

wire n2885;
// (14, 7, 'lutff_5/lout')

wire n2886;
// (11, 18, 'lutff_5/lout')

wire n2887;
// (16, 11, 'lutff_6/lout')

wire n2888;
// (15, 22, 'lutff_4/out')

wire n2889;
// (15, 22, 'lutff_4/lout')

wire n2890;
// (18, 9, 'lutff_0/lout')

wire n2891;
// (12, 19, 'lutff_7/lout')

wire n2892;
// (6, 11, 'lutff_7/lout')

wire n2893;
// (17, 23, 'lutff_1/lout')

wire n2894;
// (19, 17, 'lutff_0/out')

wire n2895;
// (22, 21, 'lutff_3/lout')

wire n2896;
// (7, 8, 'lutff_5/lout')

wire n2897;
// (21, 19, 'lutff_2/lout')

wire n2898;
// (21, 14, 'lutff_5/lout')

wire n2899;
// (12, 14, 'lutff_3/lout')

wire n2900;
// (14, 20, 'lutff_2/lout')

wire n2901;
// (10, 10, 'lutff_6/out')

wire n2902;
// (10, 10, 'lutff_6/lout')

wire n2903;
// (16, 23, 'lutff_5/lout')

wire n2904;
// (13, 20, 'lutff_2/lout')

wire n2905;
// (20, 19, 'lutff_4/lout')

wire n2906;
// (11, 12, 'lutff_7/lout')

wire n2907;
// (17, 19, 'lutff_6/out')

wire n2908;
// (17, 19, 'lutff_6/lout')

wire n2909;
// (11, 19, 'lutff_6/lout')

wire n2910;
// (16, 10, 'lutff_5/lout')

wire n2911;
// (15, 24, 'lutff_6/lout')

wire n2912;
// (12, 18, 'lutff_4/lout')

wire n2913;
// (17, 16, 'lutff_0/lout')

wire n2914;
// (19, 14, 'lutff_1/out')

wire n2915;
// (22, 20, 'lutff_0/lout')

wire n2916;
// (10, 14, 'lutff_3/lout')

wire n2917;
// (16, 24, 'lutff_1/lout')

wire n2918;
// (21, 20, 'lutff_3/lout')

wire n2919;
// (9, 17, 'lutff_5/lout')

wire n2920;
// (12, 13, 'lutff_2/lout')

wire n2921;
// (20, 12, 'lutff_2/lout')

wire n2922;
// (10, 13, 'lutff_7/lout')

wire n2923;
// (15, 11, 'lutff_0/lout')

wire n2924;
// (11, 13, 'lutff_0/lout')

wire n2925;
// (11, 16, 'lutff_7/lout')

wire n2926;
// (13, 7, 'lutff_2/out')

wire n2927;
// (15, 25, 'lutff_1/lout')

wire n2928;
// (18, 11, 'lutff_2/lout')

wire n2929;
// (15, 20, 'lutff_6/lout')

wire n2930;
// (12, 17, 'lutff_5/lout')

wire n2931;
// (17, 17, 'lutff_3/lout')

wire n2932;
// (19, 15, 'lutff_2/lout')

wire n2933;
// (22, 23, 'lutff_1/lout')

wire n2934;
// (21, 21, 'lutff_0/out')

wire n2935;
// (14, 22, 'lutff_4/lout')

wire n2936;
// (11, 9, 'lutff_5/lout')

wire n2937;
// (16, 21, 'lutff_7/lout')

wire n2938;
// (13, 22, 'lutff_0/lout')

wire n2939;
// (13, 22, 'carry_in_mux')

// Carry-In for (13 22)
assign n2939 = 0;

wire n2940;
// (15, 8, 'lutff_1/lout')

wire n2941;
// (20, 17, 'lutff_6/lout')

wire n2942;
// (23, 20, 'lutff_4/lout')

wire n2943;
// (11, 10, 'lutff_1/lout')

wire n2944;
// (9, 14, 'lutff_2/lout')

wire n2945;
// (14, 18, 'lutff_1/lout')

wire n2946;
// (17, 18, 'lutff_2/out')

wire n2947;
// (17, 18, 'lutff_2/lout')

wire n2948;
// (19, 12, 'lutff_3/lout')

wire n2949;
// (21, 22, 'lutff_1/lout')

wire n2950;
// (14, 17, 'lutff_5/lout')

wire n2951;
// (17, 12, 'lutff_1/out')

wire n2952;
// (11, 22, 'lutff_4/lout')

wire n2953;
// (10, 15, 'lutff_5/lout')

wire n2954;
// (16, 20, 'lutff_0/lout')

wire n2955;
// (21, 24, 'lutff_0/lout')

wire n2956;
// (15, 18, 'lutff_7/lout')

wire n2957;
// (18, 14, 'lutff_2/out')

wire n2958;
// (20, 16, 'lutff_1/lout')

wire n2959;
// (12, 20, 'lutff_7/lout')

wire n2960;
// (20, 13, 'lutff_6/lout')

wire n2961;
// (11, 11, 'lutff_2/lout')

wire n2962;
// (22, 18, 'lutff_3/lout')

wire n2963;
// (10, 17, 'lutff_1/lout')

wire n2964;
// (9, 15, 'lutff_5/out')

wire n2965;
// (13, 9, 'lutff_0/lout')

wire n2966;
// (21, 10, 'lutff_4/out')

wire n2967;
// (18, 13, 'lutff_4/lout')

wire n2968;
// (12, 23, 'lutff_3/out')

wire n2969;
// (12, 23, 'lutff_3/lout')

wire n2970;
// (14, 13, 'lutff_0/lout')

wire n2971;
// (19, 22, 'lutff_5/lout')

wire n2972;
// (19, 13, 'lutff_4/lout')

wire n2973;
// (16, 16, 'lutff_5/lout')

wire n2974;
// (7, 12, 'lutff_1/lout')

wire n2975;
// (15, 13, 'lutff_3/lout')

wire n2976;
// (20, 20, 'lutff_6/lout')

wire n2977;
// (14, 16, 'lutff_6/lout')

wire n2978;
// (17, 13, 'lutff_2/lout')

wire n2979;
// (16, 19, 'lutff_1/lout')

wire n2980;
// (15, 19, 'lutff_4/lout')

wire n2981;
// (18, 17, 'lutff_3/lout')

wire n2982;
// (15, 14, 'lutff_7/lout')

wire n2983;
// (20, 23, 'lutff_0/lout')

wire n2984;
// (10, 16, 'lutff_2/lout')

wire n2985;
// (13, 10, 'lutff_1/lout')

wire n2986;
// (21, 11, 'lutff_3/lout')

wire n2987;
// (18, 12, 'lutff_7/lout')

wire n2988;
// (12, 22, 'lutff_0/out')

wire n2989;
// (12, 22, 'lutff_0/lout')

wire n2990;
// (14, 12, 'lutff_3/lout')

wire n2991;
// (19, 23, 'lutff_6/lout')

wire n2992;
// (19, 10, 'lutff_5/lout')

wire n2993;
// (22, 16, 'lutff_4/lout')

wire n2994;
// (14, 19, 'lutff_7/lout')

wire n2995;
// (17, 14, 'lutff_3/out')

wire n2996;
// (19, 24, 'lutff_4/lout')

wire n2997;
// (11, 20, 'lutff_6/lout')

wire n2998;
// (16, 18, 'lutff_2/lout')

wire n2999;
// (15, 16, 'lutff_5/lout')

wire n3000;
// (15, 15, 'lutff_4/lout')

wire n3001;
// (18, 16, 'lutff_0/out')

wire n3002;
// (18, 16, 'lutff_0/lout')

wire n3003;
// (18, 16, 'carry_in_mux')

// Carry-In for (18 16)
assign n3003 = 0;

wire n3004;
// (20, 22, 'lutff_3/out')

wire n3005;
// (17, 24, 'lutff_3/out')

wire n3006;
// (17, 24, 'lutff_3/lout')

wire n3007;
// (10, 19, 'lutff_3/lout')

wire n3008;
// (13, 11, 'lutff_6/lout')

wire n3009;
// (21, 12, 'lutff_2/lout')

wire n3010;
// (18, 15, 'lutff_6/lout')

wire n3011;
// (12, 21, 'lutff_1/lout')

wire n3012;
// (19, 20, 'lutff_7/lout')

wire n3013;
// (19, 11, 'lutff_6/lout')

wire n3014;
// (22, 19, 'lutff_5/lout')

wire n3015;
// (17, 15, 'lutff_4/lout')

wire n3016;
// (16, 17, 'lutff_3/lout')

wire n3017;
// (22, 13, 'lutff_1/lout')

wire n3018;
// (15, 17, 'lutff_2/lout')

wire n3019;
// (15, 12, 'lutff_5/lout')

wire n3020;
// (18, 19, 'lutff_1/lout')

wire n3021;
// (20, 21, 'lutff_2/lout')

wire n3022;
// (17, 25, 'lutff_0/lout')

wire n3023;
// (24, 14, 'lutff_6/lout')

wire n3024;
// (21, 13, 'lutff_1/out')

wire n3025;
// (17, 11, 'lutff_1/out')

wire n3026;
// (19, 21, 'lutff_0/lout')

wire n3027;
// (11, 17, 'lutff_6/out')

wire n3028;
// (23, 14, 'lutff_4/lout')

wire n3029;
// (24, 17, 'lutff_4/lout')

wire n3030;
// (15, 21, 'lutff_7/lout')

wire n3031;
// (12, 10, 'lutff_3/lout')

wire n3032;
// (17, 8, 'lutff_5/lout')

wire n3033;
// (11, 18, 'lutff_0/lout')

wire n3034;
// (11, 18, 'carry_in_mux')

// Carry-In for (11 18)
assign n3034 = 0;

wire n3035;
// (22, 12, 'lutff_2/lout')

wire n3036;
// (13, 16, 'lutff_2/lout')

wire n3037;
// (15, 22, 'lutff_3/out')

wire n3038;
// (15, 22, 'lutff_3/lout')

wire n3039;
// (18, 9, 'lutff_7/lout')

wire n3040;
// (18, 18, 'lutff_6/out')

wire n3041;
// (6, 11, 'lutff_2/lout')

wire n3042;
// (14, 10, 'lutff_2/lout')

wire n3043;
// (19, 17, 'lutff_5/out')

wire n3044;
// (22, 21, 'lutff_6/lout')

wire n3045;
// (5, 17, 'lutff_3/lout')

wire n3046;
// (21, 14, 'lutff_0/out')

wire n3047;
// (20, 26, 'lutff_2/lout')

wire n3048;
// (14, 20, 'lutff_7/lout')

wire n3049;
// (14, 9, 'lutff_4/out')

wire n3050;
// (17, 20, 'lutff_0/lout')

wire n3051;
// (19, 18, 'lutff_1/out')

wire n3052;
// (10, 10, 'lutff_3/lout')

wire n3053;
// (23, 15, 'lutff_7/lout')

wire n3054;
// (21, 16, 'lutff_3/out')

wire n3055;
// (15, 10, 'lutff_6/lout')

wire n3056;
// (18, 22, 'lutff_3/lout')

wire n3057;
// (11, 19, 'lutff_3/lout')

wire n3058;
// (9, 12, 'lutff_7/lout')

wire n3059;
// (22, 15, 'lutff_3/lout')

wire n3060;
// (13, 17, 'lutff_1/lout')

wire n3061;
// (15, 23, 'lutff_0/lout')

wire n3062;
// (18, 21, 'lutff_7/lout')

wire n3063;
// (19, 14, 'lutff_4/out')

wire n3064;
// (22, 20, 'lutff_5/lout')

wire n3065;
// (5, 18, 'lutff_2/lout')

wire n3066;
// (16, 24, 'lutff_6/lout')

wire n3067;
// (10, 20, 'lutff_6/lout')

wire n3068;
// (20, 25, 'lutff_3/lout')

wire n3069;
// (20, 12, 'lutff_7/lout')

wire n3070;
// (19, 19, 'lutff_2/lout')

wire n3071;
// (10, 13, 'lutff_2/lout')

wire n3072;
// (23, 12, 'lutff_6/lout')

wire n3073;
// (7, 10, 'lutff_3/lout')

wire n3074;
// (21, 17, 'lutff_0/lout')

wire n3075;
// (15, 11, 'lutff_5/lout')

wire n3076;
// (18, 25, 'lutff_2/lout')

wire n3077;
// (17, 7, 'lutff_0/lout')

wire n3078;
// (20, 15, 'lutff_3/lout')

wire n3079;
// (17, 10, 'lutff_7/lout')

wire n3080;
// (22, 14, 'lutff_4/lout')

wire n3081;
// (13, 18, 'lutff_0/lout')

wire n3082;
// (13, 18, 'carry_in_mux')

// Carry-In for (13 18)
assign n3082 = 0;

wire n3083;
// (15, 20, 'lutff_1/lout')

wire n3084;
// (18, 20, 'lutff_4/lout')

wire n3085;
// (11, 14, 'lutff_1/lout')

wire n3086;
// (16, 7, 'lutff_2/lout')

wire n3087;
// (19, 15, 'lutff_7/lout')

wire n3088;
// (22, 23, 'lutff_4/lout')

wire n3089;
// (15, 26, 'lutff_0/lout')

wire n3090;
// (12, 12, 'lutff_2/lout')

wire n3091;
// (17, 22, 'lutff_2/lout')

wire n3092;
// (14, 11, 'lutff_6/lout')

wire n3093;
// (19, 16, 'lutff_3/lout')

wire n3094;
// (10, 12, 'lutff_1/lout')

wire n3095;
// (22, 10, 'lutff_1/lout')

wire n3096;
// (21, 18, 'lutff_1/lout')

wire n3097;
// (12, 15, 'lutff_4/lout')

wire n3098;
// (18, 24, 'lutff_1/lout')

wire n3099;
// (20, 14, 'lutff_0/out')

wire n3100;
// (13, 8, 'lutff_6/lout')

wire n3101;
// (13, 19, 'lutff_7/lout')

wire n3102;
// (18, 23, 'lutff_5/lout')

wire n3103;
// (14, 18, 'lutff_6/lout')

wire n3104;
// (11, 15, 'lutff_2/lout')

wire n3105;
// (14, 7, 'lutff_1/lout')

wire n3106;
// (12, 19, 'lutff_3/lout')

wire n3107;
// (14, 17, 'lutff_0/lout')

wire n3108;
// (17, 12, 'lutff_4/lout')

wire n3109;
// (17, 23, 'lutff_5/lout')

wire n3110;
// (10, 15, 'lutff_0/lout')

wire n3111;
// (10, 15, 'carry_in_mux')

// Carry-In for (10 15)
assign n3111 = 0;

wire n3112;
// (21, 19, 'lutff_6/lout')

wire n3113;
// (13, 23, 'lutff_4/out')

wire n3114;
// (13, 23, 'lutff_4/lout')

wire n3115;
// (15, 9, 'lutff_3/lout')

wire n3116;
// (12, 14, 'lutff_7/lout')

wire n3117;
// (6, 16, 'lutff_0/lout')

wire n3118;
// (20, 13, 'lutff_1/out')

wire n3119;
// (16, 23, 'lutff_1/lout')

wire n3120;
// (10, 17, 'lutff_4/lout')

wire n3121;
// (13, 20, 'lutff_6/lout')

wire n3122;
// (18, 13, 'lutff_3/out')

wire n3123;
// (20, 19, 'lutff_0/lout')

wire n3124;
// (14, 13, 'lutff_7/lout')

wire n3125;
// (11, 12, 'lutff_3/lout')

wire n3126;
// (17, 19, 'lutff_2/out')

wire n3127;
// (17, 19, 'lutff_2/lout')

wire n3128;
// (19, 13, 'lutff_1/out')

wire n3129;
// (22, 17, 'lutff_2/out')

wire n3130;
// (15, 24, 'lutff_2/lout')

wire n3131;
// (12, 18, 'lutff_0/lout')

wire n3132;
// (17, 13, 'lutff_7/lout')

wire n3133;
// (14, 16, 'lutff_3/lout')

wire n3134;
// (17, 16, 'lutff_4/out')

wire n3135;
// (7, 9, 'lutff_6/lout')

wire n3136;
// (21, 20, 'lutff_7/lout')

wire n3137;
// (13, 24, 'lutff_5/out')

wire n3138;
// (13, 24, 'lutff_5/lout')

wire n3139;
// (15, 14, 'lutff_2/lout')

wire n3140;
// (18, 17, 'lutff_6/lout')

wire n3141;
// (12, 13, 'lutff_6/lout')

wire n3142;
// (16, 22, 'lutff_2/lout')

wire n3143;
// (10, 16, 'lutff_7/lout')

wire n3144;
// (13, 10, 'lutff_4/lout')

wire n3145;
// (18, 12, 'lutff_0/lout')

wire n3146;
// (14, 12, 'lutff_4/out')

wire n3147;
// (11, 13, 'lutff_4/lout')

wire n3148;
// (19, 10, 'lutff_0/lout')

wire n3149;
// (22, 16, 'lutff_1/out')

wire n3150;
// (15, 25, 'lutff_5/lout')

wire n3151;
// (12, 17, 'lutff_1/lout')

wire n3152;
// (14, 19, 'lutff_2/lout')

wire n3153;
// (17, 14, 'lutff_6/out')

wire n3154;
// (17, 17, 'lutff_7/lout')

wire n3155;
// (21, 21, 'lutff_4/lout')

wire n3156;
// (15, 15, 'lutff_1/lout')

wire n3157;
// (11, 9, 'lutff_1/lout')

wire n3158;
// (16, 21, 'lutff_3/lout')

wire n3159;
// (10, 19, 'lutff_6/lout')

wire n3160;
// (13, 11, 'lutff_3/lout')

wire n3161;
// (13, 22, 'lutff_4/lout')

wire n3162;
// (18, 15, 'lutff_1/lout')

wire n3163;
// (20, 17, 'lutff_2/lout')

wire n3164;
// (11, 10, 'lutff_5/lout')

wire n3165;
// (19, 11, 'lutff_3/lout')

wire n3166;
// (17, 15, 'lutff_1/lout')

wire n3167;
// (19, 25, 'lutff_0/lout')

wire n3168;
// (17, 18, 'lutff_6/out')

wire n3169;
// (17, 18, 'lutff_6/lout')

wire n3170;
// (22, 13, 'lutff_4/lout')

wire n3171;
// (21, 22, 'lutff_5/lout')

wire n3172;
// (15, 12, 'lutff_0/lout')

wire n3173;
// (18, 19, 'lutff_4/lout')

wire n3174;
// (11, 22, 'lutff_0/lout')

wire n3175;
// (16, 15, 'lutff_5/lout')

wire n3176;
// (16, 20, 'lutff_4/lout')

wire n3177;
// (13, 12, 'lutff_2/lout')

wire n3178;
// (15, 18, 'lutff_3/lout')

wire n3179;
// (20, 16, 'lutff_5/lout')

wire n3180;
// (12, 20, 'lutff_3/lout')

wire n3181;
// (17, 11, 'lutff_6/lout')

wire n3182;
// (11, 11, 'lutff_6/lout')

wire n3183;
// (23, 14, 'lutff_3/lout')

wire n3184;
// (12, 23, 'lutff_7/out')

wire n3185;
// (12, 23, 'lutff_7/lout')

wire n3186;
// (19, 22, 'lutff_1/lout')

wire n3187;
// (16, 16, 'lutff_1/lout')

wire n3188;
// (22, 12, 'lutff_7/lout')

wire n3189;
// (7, 12, 'lutff_5/lout')

wire n3190;
// (18, 18, 'lutff_3/lout')

wire n3191;
// (20, 20, 'lutff_2/lout')

wire n3192;
// (14, 10, 'lutff_7/lout')

wire n3193;
// (16, 14, 'lutff_6/lout')

wire n3194;
// (5, 17, 'lutff_4/lout')

wire n3195;
// (16, 19, 'lutff_5/lout')

wire n3196;
// (15, 19, 'lutff_0/lout')

wire n3197;
// (14, 9, 'lutff_3/out')

wire n3198;
// (17, 20, 'lutff_7/lout')

wire n3199;
// (23, 15, 'lutff_0/lout')

wire n3200;
// (24, 16, 'lutff_0/lout')

wire n3201;
// (21, 16, 'lutff_6/out')

wire n3202;
// (21, 11, 'lutff_7/lout')

wire n3203;
// (12, 22, 'lutff_4/out')

wire n3204;
// (12, 22, 'lutff_4/lout')

wire n3205;
// (19, 23, 'lutff_2/lout')

wire n3206;
// (22, 15, 'lutff_6/lout')

wire n3207;
// (18, 21, 'lutff_2/lout')

wire n3208;
// (20, 11, 'lutff_3/lout')

wire n3209;
// (11, 20, 'lutff_2/lout')

wire n3210;
// (16, 13, 'lutff_7/lout')

wire n3211;
// (5, 18, 'lutff_5/lout')

wire n3212;
// (16, 18, 'lutff_6/lout')

wire n3213;
// (10, 20, 'lutff_3/lout')

wire n3214;
// (15, 16, 'lutff_1/lout')

wire n3215;
// (21, 15, 'lutff_4/lout')

wire n3216;
// (20, 25, 'lutff_6/lout')

wire n3217;
// (20, 22, 'lutff_7/lout')

wire n3218;
// (17, 24, 'lutff_7/out')

wire n3219;
// (17, 24, 'lutff_7/lout')

wire n3220;
// (23, 12, 'lutff_1/lout')

wire n3221;
// (24, 15, 'lutff_1/lout')

wire n3222;
// (7, 10, 'lutff_6/lout')

wire n3223;
// (21, 17, 'lutff_5/lout')

wire n3224;
// (21, 12, 'lutff_6/lout')

wire n3225;
// (12, 21, 'lutff_5/lout')

wire n3226;
// (17, 10, 'lutff_2/lout')

wire n3227;
// (19, 20, 'lutff_3/lout')

wire n3228;
// (22, 14, 'lutff_1/lout')

wire n3229;
// (18, 20, 'lutff_1/out')

wire n3230;
// (20, 10, 'lutff_0/lout')

wire n3231;
// (23, 16, 'lutff_7/lout')

wire n3232;
// (11, 14, 'lutff_4/lout')

wire n3233;
// (16, 12, 'lutff_0/lout')

wire n3234;
// (5, 19, 'lutff_2/lout')

wire n3235;
// (16, 17, 'lutff_7/lout')

wire n3236;
// (15, 17, 'lutff_6/lout')

wire n3237;
// (20, 24, 'lutff_1/lout')

wire n3238;
// (12, 12, 'lutff_7/lout')

wire n3239;
// (20, 21, 'lutff_6/lout')

wire n3240;
// (17, 22, 'lutff_5/lout')

wire n3241;
// (24, 14, 'lutff_2/lout')

wire n3242;
// (22, 10, 'lutff_6/lout')

wire n3243;
// (21, 18, 'lutff_4/lout')

wire n3244;
// (21, 13, 'lutff_5/out')

wire n3245;
// (12, 15, 'lutff_3/lout')

wire n3246;
// (19, 21, 'lutff_4/lout')

wire n3247;
// (10, 11, 'lutff_0/lout')

wire n3248;
// (15, 21, 'lutff_3/lout')

wire n3249;
// (18, 23, 'lutff_0/lout')

wire n3250;
// (23, 17, 'lutff_0/lout')

wire n3251;
// (11, 15, 'lutff_7/lout')

wire n3252;
// (14, 7, 'lutff_4/lout')

wire n3253;
// (11, 18, 'lutff_4/lout')

wire n3254;
// (16, 11, 'lutff_1/lout')

wire n3255;
// (15, 22, 'lutff_7/out')

wire n3256;
// (15, 22, 'lutff_7/lout')

wire n3257;
// (18, 9, 'lutff_3/lout')

wire n3258;
// (12, 19, 'lutff_6/lout')

wire n3259;
// (6, 11, 'lutff_6/lout')

wire n3260;
// (17, 23, 'lutff_2/lout')

wire n3261;
// (19, 17, 'lutff_1/out')

wire n3262;
// (22, 21, 'lutff_2/lout')

wire n3263;
// (21, 19, 'lutff_3/out')

wire n3264;
// (21, 14, 'lutff_4/lout')

wire n3265;
// (9, 16, 'lutff_1/lout')

wire n3266;
// (12, 14, 'lutff_0/lout')

wire n3267;
// (12, 14, 'carry_in_mux')

// Carry-In for (12 14)
assign n3267 = 0;

wire n3268;
// (14, 20, 'lutff_3/lout')

wire n3269;
// (19, 18, 'lutff_5/lout')

wire n3270;
// (10, 10, 'lutff_7/out')

wire n3271;
// (10, 10, 'lutff_7/lout')

wire n3272;
// (16, 23, 'lutff_4/lout')

wire n3273;
// (15, 10, 'lutff_2/lout')

wire n3274;
// (20, 19, 'lutff_7/lout')

wire n3275;
// (20, 8, 'lutff_6/lout')

wire n3276;
// (11, 12, 'lutff_6/lout')

wire n3277;
// (17, 19, 'lutff_7/out')

wire n3278;
// (17, 19, 'lutff_7/lout')

wire n3279;
// (11, 19, 'lutff_7/lout')

wire n3280;
// (16, 10, 'lutff_2/lout')

wire n3281;
// (9, 12, 'lutff_3/lout')

wire n3282;
// (15, 24, 'lutff_5/lout')

wire n3283;
// (12, 18, 'lutff_5/lout')

wire n3284;
// (17, 16, 'lutff_3/lout')

wire n3285;
// (19, 14, 'lutff_0/lout')

wire n3286;
// (22, 20, 'lutff_1/lout')

wire n3287;
// (16, 24, 'lutff_2/lout')

wire n3288;
// (21, 20, 'lutff_2/lout')

wire n3289;
// (12, 13, 'lutff_1/lout')

wire n3290;
// (14, 23, 'lutff_2/lout')

wire n3291;
// (20, 12, 'lutff_3/lout')

wire n3292;
// (19, 19, 'lutff_6/lout')

wire n3293;
// (10, 13, 'lutff_6/lout')

wire n3294;
// (15, 11, 'lutff_1/lout')

wire n3295;
// (20, 18, 'lutff_4/lout')

wire n3296;
// (20, 15, 'lutff_7/lout')

wire n3297;
// (11, 13, 'lutff_1/lout')

wire n3298;
// (11, 16, 'lutff_6/lout')

wire n3299;
// (13, 7, 'lutff_3/lout')

wire n3300;
// (15, 25, 'lutff_2/lout')

wire n3301;
// (18, 11, 'lutff_1/lout')

wire n3302;
// (15, 20, 'lutff_5/lout')

wire n3303;
// (12, 17, 'lutff_4/lout')

wire n3304;
// (17, 17, 'lutff_0/lout')

wire n3305;
// (19, 15, 'lutff_3/out')

wire n3306;
// (22, 23, 'lutff_0/lout')

wire n3307;
// (21, 21, 'lutff_1/out')

wire n3308;
// (9, 18, 'lutff_3/lout')

wire n3309;
// (14, 22, 'lutff_5/lout')

wire n3310;
// (19, 16, 'lutff_7/lout')

wire n3311;
// (16, 21, 'lutff_6/lout')

wire n3312;
// (15, 8, 'lutff_0/out')

wire n3313;
// (20, 17, 'lutff_5/lout')

wire n3314;
// (20, 14, 'lutff_4/out')

wire n3315;
// (23, 20, 'lutff_3/lout')

wire n3316;
// (14, 18, 'lutff_2/lout')

wire n3317;
// (17, 18, 'lutff_1/out')

wire n3318;
// (17, 18, 'lutff_1/lout')

wire n3319;
// (19, 12, 'lutff_2/lout')

wire n3320;
// (21, 22, 'lutff_0/lout')

wire n3321;
// (17, 12, 'lutff_0/lout')

wire n3322;
// (14, 17, 'lutff_4/out')

wire n3323;
// (11, 22, 'lutff_7/lout')

wire n3324;
// (10, 15, 'lutff_4/lout')

wire n3325;
// (16, 20, 'lutff_1/lout')

wire n3326;
// (15, 18, 'lutff_6/lout')

wire n3327;
// (13, 23, 'lutff_0/out')

wire n3328;
// (13, 23, 'lutff_0/lout')

wire n3329;
// (18, 14, 'lutff_3/lout')

wire n3330;
// (20, 16, 'lutff_2/lout')

wire n3331;
// (20, 13, 'lutff_5/lout')

wire n3332;
// (11, 11, 'lutff_3/lout')

wire n3333;
// (22, 18, 'lutff_4/out')

wire n3334;
// (10, 17, 'lutff_0/lout')

wire n3335;
// (9, 15, 'lutff_6/lout')

wire n3336;
// (18, 13, 'lutff_7/lout')

wire n3337;
// (12, 23, 'lutff_2/out')

wire n3338;
// (12, 23, 'lutff_2/lout')

wire n3339;
// (14, 13, 'lutff_3/lout')

wire n3340;
// (19, 22, 'lutff_4/lout')

wire n3341;
// (19, 13, 'lutff_5/out')

wire n3342;
// (22, 17, 'lutff_6/lout')

wire n3343;
// (16, 16, 'lutff_6/lout')

wire n3344;
// (20, 20, 'lutff_7/lout')

wire n3345;
// (14, 16, 'lutff_7/lout')

wire n3346;
// (17, 13, 'lutff_3/out')

wire n3347;
// (16, 19, 'lutff_0/lout')

wire n3348;
// (9, 11, 'lutff_3/lout')

wire n3349;
// (15, 19, 'lutff_5/lout')

wire n3350;
// (13, 24, 'lutff_1/out')

wire n3351;
// (13, 24, 'lutff_1/lout')

wire n3352;
// (18, 17, 'lutff_2/lout')

wire n3353;
// (20, 23, 'lutff_3/lout')

wire n3354;
// (10, 16, 'lutff_3/lout')

wire n3355;
// (13, 10, 'lutff_0/lout')

wire n3356;
// (18, 12, 'lutff_4/lout')

wire n3357;
// (12, 22, 'lutff_1/out')

wire n3358;
// (12, 22, 'lutff_1/lout')

wire n3359;
// (14, 12, 'lutff_0/out')

wire n3360;
// (19, 23, 'lutff_7/lout')

wire n3361;
// (19, 10, 'lutff_4/lout')

wire n3362;
// (22, 16, 'lutff_5/out')

wire n3363;
// (20, 11, 'lutff_6/lout')

wire n3364;
// (17, 14, 'lutff_2/lout')

wire n3365;
// (14, 19, 'lutff_6/lout')

wire n3366;
// (19, 24, 'lutff_3/lout')

wire n3367;
// (11, 20, 'lutff_5/lout')

wire n3368;
// (16, 18, 'lutff_3/lout')

wire n3369;
// (15, 16, 'lutff_4/lout')

wire n3370;
// (15, 15, 'lutff_5/lout')

wire n3371;
// (18, 16, 'lutff_1/lout')

wire n3372;
// (20, 22, 'lutff_0/lout')

wire n3373;
// (17, 24, 'lutff_2/out')

wire n3374;
// (17, 24, 'lutff_2/lout')

wire n3375;
// (10, 19, 'lutff_2/lout')

wire n3376;
// (18, 15, 'lutff_5/out')

wire n3377;
// (12, 21, 'lutff_0/lout')

wire n3378;
// (12, 21, 'carry_in_mux')

// Carry-In for (12 21)
assign n3378 = 0;

wire n3379;
// (14, 15, 'lutff_1/lout')

wire n3380;
// (19, 20, 'lutff_6/lout')

wire n3381;
// (19, 11, 'lutff_7/lout')

wire n3382;
// (22, 19, 'lutff_4/lout')

wire n3383;
// (24, 18, 'lutff_2/lout')

wire n3384;
// (17, 15, 'lutff_5/out')

wire n3385;
// (16, 17, 'lutff_2/lout')

wire n3386;
// (22, 13, 'lutff_0/out')

wire n3387;
// (15, 17, 'lutff_3/lout')

wire n3388;
// (15, 12, 'lutff_4/lout')

wire n3389;
// (18, 19, 'lutff_0/lout')

wire n3390;
// (20, 21, 'lutff_1/lout')

wire n3391;
// (17, 25, 'lutff_1/lout')

wire n3392;
// (16, 15, 'lutff_1/lout')

wire n3393;
// (23, 13, 'lutff_3/lout')

wire n3394;
// (24, 14, 'lutff_7/lout')

wire n3395;
// (17, 11, 'lutff_2/lout')

wire n3396;
// (19, 21, 'lutff_1/lout')

wire n3397;
// (11, 17, 'lutff_7/lout')

wire n3398;
// (23, 14, 'lutff_7/lout')

wire n3399;
// (24, 17, 'lutff_3/lout')

wire n3400;
// (17, 8, 'lutff_4/lout')

wire n3401;
// (11, 18, 'lutff_3/lout')

wire n3402;
// (22, 12, 'lutff_3/lout')

wire n3403;
// (13, 16, 'lutff_5/lout')

wire n3404;
// (15, 22, 'lutff_2/out')

wire n3405;
// (15, 22, 'lutff_2/lout')

wire n3406;
// (18, 9, 'lutff_6/lout')

wire n3407;
// (18, 18, 'lutff_7/lout')

wire n3408;
// (6, 11, 'lutff_1/lout')

wire n3409;
// (23, 18, 'lutff_1/lout')

wire n3410;
// (14, 10, 'lutff_3/lout')

wire n3411;
// (19, 17, 'lutff_6/lout')

wire n3412;
// (16, 14, 'lutff_2/lout')

wire n3413;
// (5, 17, 'lutff_0/lout')

// Carry-In for (5 17)
assign n85 = 1;

wire n3414;
// (14, 20, 'lutff_4/lout')

wire n3415;
// (17, 20, 'lutff_3/lout')

wire n3416;
// (19, 18, 'lutff_0/lout')

wire n3417;
// (23, 15, 'lutff_4/lout')

wire n3418;
// (21, 16, 'lutff_2/lout')

wire n3419;
// (18, 22, 'lutff_4/lout')

wire n3420;
// (11, 19, 'lutff_0/lout')

wire n3421;
// (22, 15, 'lutff_2/lout')

wire n3422;
// (13, 17, 'lutff_6/lout')

wire n3423;
// (18, 21, 'lutff_6/lout')

wire n3424;
// (19, 14, 'lutff_7/lout')

wire n3425;
// (16, 13, 'lutff_3/lout')

wire n3426;
// (5, 18, 'lutff_1/lout')

wire n3427;
// (10, 20, 'lutff_7/lout')

wire n3428;
// (13, 14, 'lutff_4/lout')

wire n3429;
// (21, 15, 'lutff_0/lout')

wire n3430;
// (20, 25, 'lutff_2/lout')

wire n3431;
// (17, 21, 'lutff_0/lout')

wire n3432;
// (19, 19, 'lutff_3/lout')

wire n3433;
// (23, 12, 'lutff_5/lout')

wire n3434;
// (21, 17, 'lutff_1/lout')

wire n3435;
// (18, 25, 'lutff_5/lout')

wire n3436;
// (20, 15, 'lutff_2/lout')

wire n3437;
// (11, 16, 'lutff_1/lout')

wire n3438;
// (22, 14, 'lutff_5/lout')

wire n3439;
// (13, 18, 'lutff_7/lout')

wire n3440;
// (15, 20, 'lutff_0/lout')

wire n3441;
// (15, 20, 'carry_in_mux')

// Carry-In for (15 20)
assign n3441 = 0;

wire n3442;
// (18, 20, 'lutff_5/lout')

wire n3443;
// (23, 16, 'lutff_3/lout')

wire n3444;
// (11, 14, 'lutff_0/out')

wire n3445;
// (11, 14, 'lutff_0/lout')

wire n3446;
// (11, 14, 'carry_in_mux')

// Carry-In for (11 14)
assign n3446 = 1;

wire n3447;
// (16, 7, 'lutff_5/lout')

wire n3448;
// (19, 15, 'lutff_4/lout')

wire n3449;
// (16, 12, 'lutff_4/lout')

wire n3450;
// (10, 23, 'lutff_6/lout')

wire n3451;
// (12, 12, 'lutff_3/lout')

wire n3452;
// (14, 22, 'lutff_2/lout')

wire n3453;
// (17, 22, 'lutff_1/lout')

wire n3454;
// (19, 16, 'lutff_2/lout')

wire n3455;
// (22, 10, 'lutff_2/lout')

wire n3456;
// (7, 11, 'lutff_1/lout')

wire n3457;
// (21, 18, 'lutff_0/out')

wire n3458;
// (12, 15, 'lutff_7/lout')

wire n3459;
// (18, 24, 'lutff_6/lout')

wire n3460;
// (15, 7, 'lutff_2/lout')

wire n3461;
// (20, 14, 'lutff_1/out')

wire n3462;
// (13, 19, 'lutff_0/lout')

wire n3463;
// (18, 23, 'lutff_4/lout')

wire n3464;
// (14, 18, 'lutff_7/lout')

wire n3465;
// (23, 17, 'lutff_4/lout')

wire n3466;
// (11, 15, 'lutff_3/lout')

wire n3467;
// (14, 7, 'lutff_0/lout')

wire n3468;
// (14, 7, 'carry_in_mux')

// Carry-In for (14 7)
assign n3468 = 0;

wire n3469;
// (19, 12, 'lutff_5/lout')

wire n3470;
// (16, 11, 'lutff_5/lout')

wire n3471;
// (12, 19, 'lutff_2/lout')

wire n3472;
// (17, 12, 'lutff_7/lout')

wire n3473;
// (14, 17, 'lutff_3/out')

wire n3474;
// (17, 23, 'lutff_6/lout')

wire n3475;
// (13, 23, 'lutff_5/out')

wire n3476;
// (13, 23, 'lutff_5/lout')

wire n3477;
// (12, 14, 'lutff_4/lout')

wire n3478;
// (20, 13, 'lutff_0/lout')

wire n3479;
// (16, 23, 'lutff_0/lout')

wire n3480;
// (10, 17, 'lutff_7/out')

wire n3481;
// (10, 17, 'lutff_7/lout')

wire n3482;
// (13, 20, 'lutff_1/lout')

wire n3483;
// (18, 13, 'lutff_2/out')

wire n3484;
// (20, 19, 'lutff_3/lout')

wire n3485;
// (14, 13, 'lutff_6/lout')

wire n3486;
// (23, 22, 'lutff_5/lout')

wire n3487;
// (17, 19, 'lutff_3/out')

wire n3488;
// (17, 19, 'lutff_3/lout')

wire n3489;
// (19, 13, 'lutff_2/out')

wire n3490;
// (16, 10, 'lutff_6/lout')

wire n3491;
// (15, 24, 'lutff_1/lout')

wire n3492;
// (12, 18, 'lutff_1/lout')

wire n3493;
// (14, 16, 'lutff_0/lout')

wire n3494;
// (17, 13, 'lutff_4/lout')

wire n3495;
// (21, 20, 'lutff_6/lout')

wire n3496;
// (13, 24, 'lutff_4/out')

wire n3497;
// (13, 24, 'lutff_4/lout')

wire n3498;
// (9, 17, 'lutff_6/lout')

wire n3499;
// (12, 13, 'lutff_5/lout')

wire n3500;
// (18, 26, 'lutff_0/lout')

wire n3501;
// (16, 22, 'lutff_3/lout')

wire n3502;
// (10, 16, 'lutff_4/lout')

wire n3503;
// (18, 12, 'lutff_1/lout')

wire n3504;
// (6, 13, 'lutff_3/lout')

wire n3505;
// (20, 18, 'lutff_0/lout')

wire n3506;
// (14, 12, 'lutff_5/out')

wire n3507;
// (11, 13, 'lutff_5/lout')

wire n3508;
// (15, 25, 'lutff_6/lout')

wire n3509;
// (12, 17, 'lutff_0/lout')

wire n3510;
// (12, 17, 'carry_in_mux')

// Carry-In for (12 17)
assign n3510 = 0;

wire n3511;
// (17, 14, 'lutff_5/lout')

wire n3512;
// (14, 19, 'lutff_1/lout')

wire n3513;
// (17, 17, 'lutff_4/lout')

wire n3514;
// (21, 21, 'lutff_5/lout')

wire n3515;
// (16, 21, 'lutff_2/lout')

wire n3516;
// (10, 19, 'lutff_5/lout')

wire n3517;
// (13, 22, 'lutff_3/lout')

wire n3518;
// (18, 15, 'lutff_0/lout')

wire n3519;
// (6, 12, 'lutff_0/lout')

wire n3520;
// (20, 17, 'lutff_1/lout')

wire n3521;
// (14, 15, 'lutff_4/lout')

wire n3522;
// (23, 20, 'lutff_7/lout')

wire n3523;
// (19, 11, 'lutff_0/lout')

wire n3524;
// (17, 15, 'lutff_2/lout')

wire n3525;
// (19, 25, 'lutff_1/lout')

wire n3526;
// (17, 18, 'lutff_5/out')

wire n3527;
// (17, 18, 'lutff_5/lout')

wire n3528;
// (22, 13, 'lutff_7/lout')

wire n3529;
// (11, 22, 'lutff_3/lout')

wire n3530;
// (16, 15, 'lutff_4/lout')

wire n3531;
// (16, 20, 'lutff_5/lout')

wire n3532;
// (15, 18, 'lutff_2/lout')

wire n3533;
// (20, 16, 'lutff_6/lout')

wire n3534;
// (17, 11, 'lutff_7/lout')

wire n3535;
// (11, 11, 'lutff_7/lout')

wire n3536;
// (23, 14, 'lutff_2/lout')

wire n3537;
// (22, 18, 'lutff_0/out')

wire n3538;
// (21, 10, 'lutff_7/lout')

wire n3539;
// (12, 23, 'lutff_6/out')

wire n3540;
// (12, 23, 'lutff_6/lout')

wire n3541;
// (19, 22, 'lutff_0/lout')

// Carry-In for (19 22)
assign n1510 = 1;

// plltype = 111
// (14,  0, "PLLCONFIG_7") DIVF_2
// (14,  0, "PLLCONFIG_9") DIVF_4
// (15,  0, "PLLCONFIG_2") DIVF_6
// (15,  0, "PLLCONFIG_3") DIVQ_0
// (15,  0, "PLLCONFIG_4") DIVQ_1
// (15,  0, "PLLCONFIG_6") FILTER_RANGE_0
// (16,  0, "PLLCONFIG_2") PLLOUT_SELECT_B_0
// (16,  0, "PLLCONFIG_5") PLLTYPE_0
// (18,  0, "PLLCONFIG_1") PLLTYPE_1
// (18,  0, "PLLCONFIG_3") PLLTYPE_2
// (18,  0, "PLLCONFIG_5") FEEDBACK_PATH_0
SB_PLL40_2F_CORE #(
  .FEEDBACK_PATH("SIMPLE"),
  .DELAY_ADJUSTMENT_MODE_FEEDBACK("FIXED"),
  .DELAY_ADJUSTMENT_MODE_RELATIVE("FIXED"),
  .PLLOUT_SELECT_PORTA("GENCLK"),
  .PLLOUT_SELECT_PORTB("GENCLK_HALF"),
  .SHIFTREG_DIV_MODE(1'b0),
  .FDA_FEEDBACK(4'b0000),
  .FDA_RELATIVE(4'b0000),
  .DIVR(4'b0000),
  .DIVF(7'b1010100),
  .DIVQ(3'b011),
  .FILTER_RANGE(3'b001),
  .ENABLE_ICEGATE_PORTA(1'b0),
  .ENABLE_ICEGATE_PORTB(1'b0),
  .TEST_MODE(1'b0)
) PLL_16_0 (
  .REFERENCECLK(io_0_16_1),
  .PLLOUTCOREA(n3),
  .PLLOUTCOREB(n1),
  .EXTFEEDBACK(1'b0),
  .DYNAMICDELAY({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
  .LOCK(n1772),
  .BYPASS(1'b0),
  .RESETB(io_0_25_1),
  .LATCHINPUTVALUE(1'b0),
  .SDO(n1773),
  .SDI(1'b0),
  .SCLK(1'b0)
);

// IO Cell (33, 14, 1)
// PAD     = io_33_14_1
// D_IN_0  = n1382
// D_IN_1  = 
// D_OUT_0 = n1017
// D_OUT_1 = 0
// OUT_ENB = n1377
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1382 = io_33_14_1;
assign io_33_14_1 = n1377 ? n1017 : 1'bz;

// IO Cell (33, 2, 1)
// PAD     = io_33_2_1
// D_IN_0  = n331
// D_IN_1  = 
// D_OUT_0 = n1016
// D_OUT_1 = 0
// OUT_ENB = n1376
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n331 = io_33_2_1;
assign io_33_2_1 = n1376 ? n1016 : 1'bz;

// IO Cell (33, 6, 1)
// PAD     = io_33_6_1
// D_IN_0  = n383
// D_IN_1  = 
// D_OUT_0 = n192
// D_OUT_1 = 0
// OUT_ENB = n1260
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n383 = io_33_6_1;
assign io_33_6_1 = n1260 ? n192 : 1'bz;

// IO Cell (31, 33, 1)
// PAD     = io_31_33_1
// D_IN_0  = n1494
// D_IN_1  = 
// D_OUT_0 = n1697
// D_OUT_1 = 0
// OUT_ENB = n1379
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1494 = io_31_33_1;
assign io_31_33_1 = n1379 ? n1697 : 1'bz;

// IO Cell (31, 33, 0)
// PAD     = io_31_33_0
// D_IN_0  = n1502
// D_IN_1  = 
// D_OUT_0 = n274
// D_OUT_1 = 0
// OUT_ENB = n1400
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1502 = io_31_33_0;
assign io_31_33_0 = n1400 ? n274 : 1'bz;

// IO Cell (33, 15, 1)
// PAD     = io_33_15_1
// D_IN_0  = n1349
// D_IN_1  = 
// D_OUT_0 = n1019
// D_OUT_1 = 0
// OUT_ENB = n1148
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1349 = io_33_15_1;
assign io_33_15_1 = n1148 ? n1019 : 1'bz;

// IO Cell (29, 33, 1)
// PAD     = io_29_33_1
// D_IN_0  = n1146
// D_IN_1  = 
// D_OUT_0 = n1022
// D_OUT_1 = 0
// OUT_ENB = n1403
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1146 = io_29_33_1;
assign io_29_33_1 = n1403 ? n1022 : 1'bz;

// IO Cell (33, 15, 0)
// PAD     = io_33_15_0
// D_IN_0  = n1388
// D_IN_1  = 
// D_OUT_0 = n1018
// D_OUT_1 = 0
// OUT_ENB = n1259
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1388 = io_33_15_0;
assign io_33_15_0 = n1259 ? n1018 : 1'bz;

// IO Cell (33, 16, 0)
// PAD     = io_33_16_0
// D_IN_0  = n1398
// D_IN_1  = 
// D_OUT_0 = n1020
// D_OUT_1 = 0
// OUT_ENB = n1402
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1398 = io_33_16_0;
assign io_33_16_0 = n1402 ? n1020 : 1'bz;

// IO Cell (29, 33, 0)
// PAD     = io_29_33_0
// D_IN_0  = n1261
// D_IN_1  = 
// D_OUT_0 = n104
// D_OUT_1 = 0
// OUT_ENB = n1380
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1261 = io_29_33_0;
assign io_29_33_0 = n1380 ? n104 : 1'bz;

// IO Cell (33, 16, 1)
// PAD     = io_33_16_1
// D_IN_0  = n1397
// D_IN_1  = 
// D_OUT_0 = n132
// D_OUT_1 = 0
// OUT_ENB = n729
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1397 = io_33_16_1;
assign io_33_16_1 = n729 ? n132 : 1'bz;

// IO Cell (30, 33, 0)
// PAD     = io_30_33_0
// D_IN_0  = n1242
// D_IN_1  = 
// D_OUT_0 = n543
// D_OUT_1 = 0
// OUT_ENB = n1378
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1242 = io_30_33_0;
assign io_30_33_0 = n1378 ? n543 : 1'bz;

// IO Cell (30, 33, 1)
// PAD     = io_30_33_1
// D_IN_0  = n1381
// D_IN_1  = 
// D_OUT_0 = n1023
// D_OUT_1 = 0
// OUT_ENB = n1024
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1381 = io_30_33_1;
assign io_30_33_1 = n1024 ? n1023 : 1'bz;

// IO Cell (33, 10, 1)
// PAD     = io_33_10_1
// D_IN_0  = n880
// D_IN_1  = 
// D_OUT_0 = n146
// D_OUT_1 = 0
// OUT_ENB = n1401
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n880 = io_33_10_1;
assign io_33_10_1 = n1401 ? n146 : 1'bz;

// IO Cell (27, 33, 0)
// PAD     = io_27_33_0
// D_IN_0  = n1011
// D_IN_1  = 
// D_OUT_0 = n1014
// D_OUT_1 = 0
// OUT_ENB = n1021
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1011 = io_27_33_0;
assign io_27_33_0 = n1021 ? n1014 : 1'bz;

// IO Cell (28, 33, 1)
// PAD     = io_28_33_1
// D_IN_0  = n1500
// D_IN_1  = 
// D_OUT_0 = n1015
// D_OUT_1 = 0
// OUT_ENB = n1404
// CLK_EN  = 1
// IN_CLK  = 0
// OUT_CLK = 0
// LATCH   = 0
// TYPE    = 100101 (LSB:MSB)
assign n1500 = io_28_33_1;
assign io_28_33_1 = n1404 ? n1015 : 1'bz;

assign n1953 = 1'b0;
assign n1967 = 1'b0;
assign n1998 = 1'b0;
assign n2012 = 1'b0;
assign n2061 = 1'b0;
assign n2068 = 1'b0;
assign n2090 = 1'b0;
assign n2202 = 1'b0;
assign n2209 = 1'b0;
assign n2215 = 1'b0;
assign n2227 = 1'b0;
assign n2258 = 1'b0;
assign n2275 = 1'b0;
assign n2291 = 1'b0;
assign n2308 = 1'b0;
assign n2338 = 1'b0;
assign n2406 = 1'b0;
assign n2419 = 1'b0;
assign n2429 = 1'b0;
assign n2464 = 1'b0;
assign n2474 = 1'b0;
assign n2492 = 1'b0;
assign n2507 = 1'b0;
assign n2538 = 1'b0;
assign n2545 = 1'b0;
assign n2550 = 1'b0;
assign n2557 = 1'b0;
assign n2568 = 1'b0;
assign n2592 = 1'b0;
assign n2607 = 1'b0;
assign n2623 = 1'b0;
assign n2637 = 1'b0;
assign n2669 = 1'b0;
assign n2724 = 1'b0;
assign n2743 = 1'b0;
assign n2755 = 1'b0;
assign n2767 = 1'b0;
assign n2797 = 1'b0;
assign n32   = 1'b1;
assign n2816 = 1'b0;
assign n2836 = 1'b0;
assign n2852 = 1'b0;
assign n2888 = 1'b0;
assign n2901 = 1'b0;
assign n2907 = 1'b0;
assign n2946 = 1'b0;
assign n2968 = 1'b0;
assign n2988 = 1'b0;
assign n3001 = 1'b0;
assign n3005 = 1'b0;
assign n3037 = 1'b0;
assign n3113 = 1'b0;
assign n3126 = 1'b0;
assign n3137 = 1'b0;
assign n3168 = 1'b0;
assign n3184 = 1'b0;
assign n3203 = 1'b0;
assign n3218 = 1'b0;
assign n3255 = 1'b0;
assign n3270 = 1'b0;
assign n3277 = 1'b0;
assign n3317 = 1'b0;
assign n3327 = 1'b0;
assign n3337 = 1'b0;
assign n3350 = 1'b0;
assign n3357 = 1'b0;
assign n3373 = 1'b0;
assign n3404 = 1'b0;
assign n3444 = 1'b0;
assign n3475 = 1'b0;
assign n3480 = 1'b0;
assign n3487 = 1'b0;
assign n3496 = 1'b0;
assign n3526 = 1'b0;
assign n3539 = 1'b0;
assign n1940 = /* LUT   16 16  2 */ n44 ? 1'b1 : 1'b0;
assign n1941 = /* LUT   22 12  4 */ n35 ? 1'b1 : 1'b0;
assign n945  = /* LUT   15 13  0 */ n778 ? n943 ? 1'b0 : n244 ? 1'b1 : 1'b0 : n943 ? n244 ? 1'b1 : 1'b0 : 1'b0;
assign n1943 = /* LUT   20 20  3 */ n42 ? 1'b1 : 1'b0;
assign n1944 = /* LUT   16 14  7 */ n59 ? n244 ? n525 ? 1'b0 : n948 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n1945 = /* LUT    5 17  5 */ n90 ? n49 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n49 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n1946 = /* LUT   16 19  4 */ n140 ? 1'b1 : 1'b0;
assign n1947 = /* LUT   15 19  1 */ n212 ? 1'b1 : 1'b0;
assign n1948 = /* LUT   17 20  6 */ n190 ? 1'b0 : 1'b1;
assign n1949 = /* LUT   23 15  1 */ n212 ? 1'b1 : 1'b0;
assign n1950 = /* LUT   24 16  1 */ n158 ? 1'b1 : 1'b0;
assign n1951 = /* LUT    7 16  7 */ io_0_20_0 ? 1'b1 : io_25_0_0 ? 1'b1 : io_0_16_0 ? 1'b1 : 1'b0;
assign n1952 = /* LUT   21 11  0 */ n159 ? 1'b1 : 1'b0;
assign n1955 = /* LUT   19 23  3 */ n272 ? n1401 ? io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0;
assign n1956 = /* LUT   10  9  5 */ n199 ? n152 ? n150 ? 1'b0 : 1'b1 : n150 ? n279 ? 1'b0 : 1'b1 : 1'b0 : n152 ? n150 ? n279 ? 1'b0 : 1'b1 : 1'b1 : 1'b0;
assign n1957 = /* LUT   22 15  5 */ n59 ? 1'b0 : n525 ? 1'b0 : n244 ? 1'b0 : n590 ? 1'b1 : 1'b0;
assign n1958 = /* LUT   20 11  2 */ n42 ? 1'b1 : 1'b0;
assign n1959 = /* LUT   19 24  7 */ n1532 ? n797 ? 1'b0 : n1501 ? 1'b0 : 1'b1 : n797 ? n1501 ? 1'b0 : 1'b1 : 1'b0;
assign n1960 = /* LUT   11 20  1 */ n248 ? 1'b0 : 1'b1;
assign n1079 = /* LUT   16 13  6 */ n59 ? 1'b1 : n440 ? n180 ? 1'b0 : 1'b1 : 1'b1;
assign n1961 = /* LUT    5 18  4 */ n97 ? n56 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n56 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n1962 = /* LUT   16 18  7 */ n218 ? 1'b1 : 1'b0;
assign n1963 = /* LUT   10 20  0 */ n44 ? 1'b1 : 1'b0;
assign n1964 = /* LUT   21 15  5 */ n42 ? 1'b1 : 1'b0;
assign n1965 = /* LUT   20 22  4 */ n1503 ? 1'b1 : n1619 ? 1'b1 : n1390 ? 1'b1 : n1391 ? 1'b1 : 1'b0;
assign n1966 = /* LUT   17 21  5 */ n724 ? n1257 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1257 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n1969 = /* LUT   23 12  0 */ n159 ? 1'b1 : 1'b0;
assign n1970 = /* LUT   24 15  0 */ n159 ? 1'b1 : 1'b0;
assign n1971 = /* LUT   21 12  1 */ n212 ? 1'b1 : 1'b0;
assign n1972 = /* LUT   12 21  4 */ n31 ? 1'b0 : 1'b1;
assign n1973 = /* LUT   17 10  1 */ 1'b0 ? 1'b1 : 1'b0;
assign n1974 = /* LUT   19 20  2 */ n1025 ? io_0_25_1 ? n1378 ? 1'b1 : n272 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n1975 = /* LUT   22 14  2 */ n44 ? 1'b1 : 1'b0;
assign n1976 = /* LUT   23 16  6 */ n140 ? 1'b1 : 1'b0;
assign n1977 = /* LUT   11 14  7 */ n457 ? n438 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n438 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n1978 = /* LUT   16 12  1 */ n770 ? 1'b0 : n212 ? 1'b1 : 1'b0;
assign n1979 = /* LUT   16 17  6 */ n140 ? 1'b1 : 1'b0;
assign n1980 = /* LUT   13 15  0 */ n579 ? 1'b1 : 1'b0;
assign n1981 = /* LUT   15 17  7 */ n218 ? 1'b1 : 1'b0;
assign n1982 = /* LUT   20 24  2 */ n1407 ? n1521 ? n1408 ? n1520 ? 1'b1 : 1'b0 : 1'b0 : n1408 ? 1'b0 : n1520 ? 1'b1 : 1'b0 : n1521 ? n1408 ? n1520 ? 1'b0 : 1'b1 : 1'b0 : n1408 ? 1'b0 : n1520 ? 1'b0 : 1'b1;
assign n1983 = /* LUT   20 21  5 */ n158 ? 1'b1 : 1'b0;
assign n1984 = /* LUT   17 22  4 */ n982 ? 1'b0 : 1'b1;
assign n1985 = /* LUT   24 14  3 */ n42 ? 1'b1 : 1'b0;
assign n1986 = /* LUT   22 10  7 */ n1707 ? n1540 ? 1'b0 : 1'b1 : n1540 ? n1537 ? 1'b0 : 1'b1 : 1'b0;
assign n1644 = /* LUT   21 13  2 */ n684 ? n1643 ? 1'b1 : n575 ? 1'b1 : 1'b0 : n1643 ? n575 ? 1'b0 : 1'b1 : 1'b0;
assign n1988 = /* LUT   12 15  2 */ n486 ? 1'b0 : 1'b1;
assign n1989 = /* LUT   19 21  5 */ n641 ? n1381 ? n1025 ? 1'b0 : 1'b1 : 1'b0 : n1349 ? n1025 ? 1'b0 : 1'b1 : 1'b0;
assign n496  = /* LUT   11 17  3 */ n494 ? 1'b0 : n246 ? n495 ? 1'b0 : n345 ? 1'b0 : 1'b1 : 1'b0;
assign n1990 = /* LUT   16  8  6 */ 1'b0 ? 1'b1 : 1'b0;
assign n1991 = /* LUT   24 17  7 */ n218 ? 1'b1 : 1'b0;
assign n1992 = /* LUT   15 21  4 */ n1000 ? 1'b0 : 1'b1;
assign n1745 = /* LUT   23 17  1 */ n1719 ? n1716 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1716 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n1994 = /* LUT   11 15  4 */ n477 ? n299 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n299 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n1995 = /* LUT   11 18  7 */ n510 ? 1'b0 : 1'b1;
assign n1996 = /* LUT   16 11  0 */ n159 ? 1'b1 : 1'b0;
assign n1997 = /* LUT   13 16  1 */ n42 ? 1'b1 : 1'b0;
assign n2000 = /* LUT   18  9  2 */ n1288 ? 1'b1 : 1'b0;
assign n2001 = /* LUT    6 11  5 */ n117 ? n72 ? 1'b0 : n81 ? 1'b0 : 1'b1 : n72 ? n81 ? 1'b0 : 1'b1 : 1'b0;
assign n2002 = /* LUT   12 24  0 */ n642 ? 1'b1 : 1'b0;
assign n2003 = /* LUT   17 23  3 */ n987 ? 1'b0 : 1'b1;
assign n2004 = /* LUT   19 17  2 */ n712 ? n1477 ? 1'b1 : 1'b0 : n502 ? 1'b1 : 1'b0;
assign n2005 = /* LUT   22 21  5 */ n158 ? 1'b1 : 1'b0;
assign n2006 = /* LUT   24 13  2 */ n218 ? 1'b1 : 1'b0;
assign n1649 = /* LUT   21 14  3 */ n1561 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1633 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1633 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2008 = /* LUT    9 16  0 */ n232 ? n234 ? n233 ? n231 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2009 = /* LUT   12 14  1 */ n469 ? 1'b0 : 1'b1;
assign n2010 = /* LUT   14 20  0 */ n852 ? n398 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n398 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n1489 = /* LUT   19 18  4 */ n966 ? n1488 ? n575 ? 1'b1 : 1'b0 : n789 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1488 ? 1'b0 : n789 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2015 = /* LUT   16 23  7 */ io_7_33_1 ? 1'b1 : 1'b0;
assign n2016 = /* LUT   15 10  5 */ n41 ? 1'b0 : n672 ? 1'b1 : n754 ? n752 ? 1'b0 : 1'b1 : 1'b0;
assign n2017 = /* LUT   20 19  6 */ n140 ? 1'b1 : 1'b0;
assign n2018 = /* LUT   18 22  0 */ n1025 ? io_0_25_1 ? n272 ? 1'b0 : 1'b1 : 1'b0 : n697 ? io_0_25_1 ? 1'b1 : 1'b0 : 1'b0;
assign n2019 = /* LUT   11 12  5 */ n429 ? 1'b1 : 1'b0;
assign n2020 = /* LUT   11 19  4 */ n261 ? 1'b0 : 1'b1;
assign n2021 = /* LUT   16 10  3 */ n1054 ? 1'b1 : 1'b0;
assign n205  = /* LUT    9 12  2 */ n80 ? n75 ? 1'b1 : n108 ? n109 ? 1'b0 : 1'b1 : 1'b0 : n108 ? n109 ? 1'b0 : 1'b1 : 1'b0;
assign n2023 = /* LUT   15 24  4 */ n1030 ? n888 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n888 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n710  = /* LUT   13 17  2 */ n269 ? 1'b0 : n514 ? 1'b0 : n268 ? 1'b0 : n516 ? 1'b0 : 1'b1;
assign n1212 = /* LUT   17 16  2 */ n1111 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1209 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1209 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n1451 = /* LUT   19 14  3 */ n792 ? n1180 ? n575 ? 1'b0 : n1095 ? 1'b0 : 1'b1 : n575 ? 1'b1 : 1'b0 : n1180 ? n575 ? 1'b0 : n1095 ? 1'b0 : 1'b1 : 1'b1;
assign n2027 = /* LUT   22 20  6 */ n1694 ? n1509 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1509 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2028 = /* LUT   16 24  3 */ io_5_33_0 ? 1'b1 : 1'b0;
assign n2029 = /* LUT   12 13  0 */ n159 ? 1'b1 : 1'b0;
assign n2030 = /* LUT   20 12  4 */ n35 ? 1'b1 : 1'b0;
assign n2031 = /* LUT   10 13  1 */ n306 ? n206 ? 1'b0 : n120 ? 1'b0 : 1'b1 : n206 ? n120 ? 1'b0 : 1'b1 : 1'b0;
assign n2032 = /* LUT   16 22  4 */ n272 ? 1'b0 : n1127 ? io_0_25_1 ? n731 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2033 = /* LUT   15 11  6 */ n921 ? 1'b1 : 1'b0;
assign n2034 = /* LUT   20 18  5 */ n1482 ? n575 ? n1600 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n1600 ? 1'b1 : 1'b0 : 1'b0;
assign n2035 = /* LUT   20 15  6 */ n1302 ? n244 ? 1'b0 : n180 ? 1'b0 : n590 ? 1'b1 : 1'b0 : 1'b0;
assign n2036 = /* LUT   11 13  2 */ n35 ? 1'b1 : 1'b0;
assign n2037 = /* LUT   11 16  5 */ n51 ? n343 ? 1'b1 : n358 ? 1'b0 : 1'b1 : n343 ? n168 ? 1'b1 : 1'b0 : n168 ? n358 ? 1'b0 : 1'b1 : 1'b0;
assign n2038 = /* LUT    9 13  1 */ n36 ? 1'b1 : 1'b0;
assign n2039 = /* LUT   15 25  3 */ n1038 ? n895 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n895 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2040 = /* LUT   13 18  3 */ n494 ? 1'b0 : 1'b1;
assign n2041 = /* LUT   18 11  0 */ n159 ? 1'b1 : 1'b0;
assign n2042 = /* LUT   15 20  4 */ n839 ? 1'b0 : 1'b1;
assign n1220 = /* LUT   17 17  1 */ n913 ? n1177 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1177 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2044 = /* LUT   16  7  1 */ n1048 ? n901 ? 1'b0 : n737 ? 1'b0 : 1'b1 : n901 ? n737 ? 1'b0 : 1'b1 : 1'b0;
assign n2045 = /* LUT   19 15  0 */ n159 ? 1'b1 : 1'b0;
assign n2046 = /* LUT   22 23  7 */ n218 ? 1'b1 : 1'b0;
assign n2047 = /* LUT    9 18  2 */ n140 ? 1'b1 : 1'b0;
assign n2048 = /* LUT   11  9  7 */ n198 ? n408 ? n151 ? n150 ? 1'b0 : 1'b1 : 1'b0 : n151 ? n150 ? 1'b0 : 1'b1 : n150 ? 1'b1 : 1'b0 : n408 ? n151 ? n150 ? 1'b0 : 1'b1 : 1'b0 : n151 ? 1'b1 : 1'b0;
assign n2049 = /* LUT   19 16  6 */ n140 ? 1'b1 : 1'b0;
assign n2050 = /* LUT   16 21  5 */ n218 ? 1'b1 : 1'b0;
assign n2051 = /* LUT   15  8  7 */ n648 ? n910 ? 1'b1 : 1'b0 : n747 ? 1'b1 : 1'b0;
assign n2052 = /* LUT    6 12  5 */ n64 ? 1'b1 : n123 ? n79 ? 1'b1 : 1'b0 : n77 ? n79 ? 1'b1 : 1'b0 : 1'b0;
assign n2053 = /* LUT   15  7  6 */ n648 ? n908 ? n647 ? 1'b0 : io_33_1_1 ? 1'b0 : 1'b1 : io_33_1_1 ? 1'b0 : 1'b1 : io_33_1_1 ? 1'b0 : 1'b1;
assign n2054 = /* LUT   18 24  2 */ n1162 ? n1412 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1412 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2055 = /* LUT   20 17  4 */ n1472 ? n1360 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1360 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2056 = /* LUT   20 14  5 */ n595 ? n705 ? n1566 ? 1'b0 : 1'b1 : 1'b0 : n1570 ? n705 ? 1'b0 : 1'b1 : 1'b1;
assign n2057 = /* LUT   23 20  2 */ n44 ? 1'b1 : 1'b0;
assign n2058 = /* LUT   11 10  3 */ n283 ? n413 ? n294 ? 1'b0 : n286 ? 1'b0 : 1'b1 : 1'b0 : n413 ? n286 ? 1'b0 : 1'b1 : 1'b0;
assign n2059 = /* LUT   13 19  4 */ n187 ? 1'b0 : 1'b1;
assign n2060 = /* LUT   14 18  3 */ n830 ? n494 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n494 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2064 = /* LUT   19 12  1 */ n590 ? n244 ? n525 ? 1'b0 : n59 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2065 = /* LUT   17 12  3 */ n756 ? n1181 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1181 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2066 = /* LUT   10 15  3 */ n334 ? n222 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n222 ? 1'b1 : 1'b0;
assign n2067 = /* LUT   16 20  2 */ n937 ? 1'b0 : n244 ? n238 ? 1'b1 : 1'b0 : 1'b0;
assign n2070 = /* LUT   15  9  0 */ n916 ? 1'b1 : 1'b0;
assign n1326 = /* LUT   18 14  4 */ n1094 ? n709 ? n930 ? 1'b0 : 1'b1 : n930 ? 1'b0 : n1236 ? 1'b0 : 1'b1 : n709 ? n930 ? 1'b0 : 1'b1 : n930 ? 1'b1 : n1236 ? 1'b0 : 1'b1;
assign n2072 = /* LUT   20 16  3 */ n42 ? 1'b1 : 1'b0;
assign n2073 = /* LUT   20 13  4 */ n1440 ? n1558 ? n930 ? 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? 1'b0 : 1'b1 : n1558 ? n930 ? n709 ? 1'b1 : 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? n709 ? 1'b1 : 1'b0 : 1'b1;
assign n2074 = /* LUT   11 11  0 */ n415 ? n285 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n285 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n1739 = /* LUT   22 18  5 */ n1586 ? n1738 ? n709 ? 1'b1 : 1'b0 : n1609 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1738 ? 1'b0 : n1609 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n2076 = /* LUT   10 17  3 */ n362 ? n243 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n243 ? 1'b1 : 1'b0;
assign n2077 = /* LUT    9 15  7 */ n225 ? n229 ? n226 ? n224 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2078 = /* LUT   13 20  5 */ n396 ? 1'b0 : 1'b1;
assign n1315 = /* LUT   18 13  6 */ n1064 ? n709 ? n930 ? 1'b0 : 1'b1 : n1074 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1074 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2080 = /* LUT   14 13  2 */ n44 ? 1'b1 : 1'b0;
assign n2081 = /* LUT   19 22  7 */ n1517 ? n1396 ? 1'b0 : n1258 ? 1'b0 : 1'b1 : n1396 ? n1258 ? 1'b0 : 1'b1 : 1'b0;
assign n2082 = /* LUT   19 13  6 */ n1303 ? n1445 ? n575 ? 1'b1 : 1'b0 : n1442 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1445 ? 1'b0 : n1442 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2083 = /* LUT   23 11  1 */ n35 ? 1'b1 : 1'b0;
assign n2084 = /* LUT   22 17  1 */ n712 ? n1730 ? 1'b1 : 1'b0 : n1709 ? 1'b1 : 1'b0;
assign n2085 = /* LUT   16 16  7 */ n218 ? 1'b1 : 1'b0;
assign n2086 = /* LUT   15 13  5 */ n244 ? n947 ? 1'b1 : 1'b0 : 1'b1;
assign n2087 = /* LUT   17 13  0 */ n140 ? 1'b1 : 1'b0;
assign n807  = /* LUT   14 16  4 */ n547 ? n701 ? 1'b0 : 1'b1 : 1'b0;
assign n2089 = /* LUT   16 19  3 */ n158 ? 1'b1 : 1'b0;
assign n956  = /* LUT   15 14  1 */ n540 ? n955 ? n525 ? n935 ? 1'b1 : 1'b0 : 1'b1 : n935 ? 1'b1 : 1'b0 : n955 ? n525 ? 1'b0 : 1'b1 : 1'b0;
assign n1354 = /* LUT   18 17  5 */ n1218 ? n1353 ? n930 ? 1'b0 : n709 ? 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n1353 ? n930 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n930 ? n709 ? 1'b0 : 1'b1 : 1'b1;
assign n2093 = /* LUT   20 23  2 */ n159 ? 1'b1 : 1'b0;
assign n2094 = /* LUT   10 16  0 */ n339 ? n229 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n229 ? 1'b1 : 1'b0;
assign n2095 = /* LUT   13 10  7 */ n664 ? 1'b1 : 1'b0;
assign n2096 = /* LUT   18 12  5 */ n158 ? 1'b1 : 1'b0;
assign n2097 = /* LUT   14 12  1 */ n676 ? n772 ? 1'b1 : n151 ? 1'b0 : 1'b1 : n772 ? n151 ? 1'b1 : 1'b0 : 1'b0;
assign n2098 = /* LUT   19 23  4 */ n1025 ? io_0_25_1 ? n272 ? n1402 ? 1'b1 : 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2099 = /* LUT   19 10  7 */ n218 ? 1'b1 : 1'b0;
assign n2100 = /* LUT   22 16  2 */ n1659 ? n1722 ? n575 ? 1'b1 : 1'b0 : n1467 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1722 ? 1'b0 : n1467 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2101 = /* LUT   26 17  2 */ 1'b0 ? 1'b1 : 1'b0;
assign n2102 = /* LUT   14 19  5 */ n849 ? n515 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n515 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2103 = /* LUT   17 14  1 */ n961 ? n1196 ? n575 ? 1'b1 : 1'b0 : n575 ? n714 ? 1'b1 : 1'b0 : 1'b1 : n1196 ? 1'b0 : n575 ? n714 ? 1'b1 : 1'b0 : 1'b1;
assign n2104 = /* LUT   19 24  2 */ n1527 ? n1407 ? 1'b0 : n1501 ? 1'b0 : 1'b1 : n1407 ? n1501 ? 1'b0 : 1'b1 : 1'b0;
assign n2105 = /* LUT   11 20  4 */ n251 ? 1'b0 : 1'b1;
assign n2106 = /* LUT   16 18  0 */ n159 ? 1'b1 : 1'b0;
assign n2107 = /* LUT   15 15  2 */ n44 ? 1'b1 : 1'b0;
assign n1618 = /* LUT   20 22  1 */ n697 ? n1273 ? 1'b1 : 1'b0 : 1'b1;
assign n2109 = /* LUT   10 19  1 */ n212 ? 1'b1 : 1'b0;
assign n674  = /* LUT   13 11  0 */ n568 ? 1'b0 : n562 ? n560 ? n567 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2110 = /* LUT   13 22  7 */ n271 ? 1'b0 : 1'b1;
assign n1334 = /* LUT   18 15  4 */ n1170 ? n1180 ? n1332 ? 1'b1 : 1'b0 : 1'b1 : n1180 ? n1332 ? 1'b1 : 1'b0 : 1'b0;
assign n2112 = /* LUT   14 15  0 */ n796 ? n694 ? n797 ? n693 ? 1'b1 : 1'b0 : 1'b0 : n797 ? 1'b0 : n693 ? 1'b1 : 1'b0 : n694 ? n797 ? n693 ? 1'b0 : 1'b1 : 1'b0 : n797 ? 1'b0 : n693 ? 1'b0 : 1'b1;
assign n2113 = /* LUT   19 11  4 */ n35 ? 1'b1 : 1'b0;
assign n2114 = /* LUT   22 19  3 */ n158 ? 1'b1 : 1'b0;
assign n2115 = /* LUT   17 15  6 */ n969 ? n1207 ? n575 ? 1'b1 : 1'b0 : n808 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1207 ? 1'b0 : n808 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2116 = /* LUT   11 21  3 */ n540 ? n244 ? 1'b0 : n59 ? 1'b0 : n525 ? 1'b0 : 1'b1 : 1'b0;
assign n2117 = /* LUT   16 17  1 */ n212 ? 1'b1 : 1'b0;
assign n1714 = /* LUT   22 13  3 */ n1641 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1636 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1636 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2119 = /* LUT    6  8  1 */ io_0_6_0 ? io_0_12_1 ? 1'b0 : 1'b1 : 1'b0;
assign n2120 = /* LUT   20 21  0 */ n1496 ? n1506 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1506 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n1097 = /* LUT   16 15  0 */ n778 ? n943 ? 1'b0 : n780 ? 1'b1 : 1'b0 : 1'b0;
assign n2121 = /* LUT   23 13  4 */ n1711 ? n1742 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1742 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2122 = /* LUT   24 14  4 */ n35 ? 1'b1 : 1'b0;
assign n2123 = /* LUT   13 12  1 */ n678 ? 1'b1 : 1'b0;
assign n2124 = /* LUT   14 21  6 */ n44 ? 1'b1 : 1'b0;
assign n2125 = /* LUT   12 20  0 */ n159 ? 1'b1 : 1'b0;
assign n1169 = /* LUT   17 11  3 */ n1062 ? n575 ? n430 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n430 ? 1'b1 : 1'b0 : 1'b0;
assign n2127 = /* LUT   19 21  2 */ n1025 ? 1'b0 : n1261 ? n641 ? 1'b1 : n331 ? 1'b1 : 1'b0 : n641 ? 1'b0 : n331 ? 1'b1 : 1'b0;
assign n2128 = /* LUT   23 14  6 */ n140 ? 1'b1 : 1'b0;
assign n2129 = /* LUT   24 17  2 */ n44 ? 1'b1 : 1'b0;
assign n2130 = /* LUT   21 10  3 */ n1622 ? n1627 ? 1'b0 : n1538 ? 1'b0 : n1626 ? 1'b0 : 1'b1 : 1'b0;
assign n555  = /* LUT   12 10  1 */ n152 ? n550 ? 1'b1 : 1'b0 : n551 ? 1'b1 : 1'b0;
assign n2132 = /* LUT   11 18  2 */ n505 ? 1'b0 : 1'b1;
assign n2133 = /* LUT   22 12  0 */ n159 ? 1'b1 : 1'b0;
assign n2134 = /* LUT   13 16  4 */ n140 ? 1'b1 : 1'b0;
assign n2135 = /* LUT   18 18  0 */ n1116 ? n575 ? n822 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n822 ? 1'b1 : 1'b0 : 1'b0;
assign n2136 = /* LUT    6 11  0 */ n112 ? n67 ? n81 ? 1'b1 : 1'b0 : 1'b1 : n67 ? 1'b1 : n81 ? 1'b1 : 1'b0;
assign n2137 = /* LUT   23 18  0 */ n159 ? 1'b1 : 1'b0;
assign n2138 = /* LUT   14 10  4 */ n757 ? 1'b1 : 1'b0;
assign n2139 = /* LUT   16 14  3 */ n770 ? 1'b0 : n158 ? 1'b1 : 1'b0;
assign n2140 = /* LUT    5 17  1 */ n86 ? n46 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n46 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2141 = /* LUT   13 13  2 */ n14 ? n546 ? 1'b0 : 1'b1 : 1'b0;
assign n2142 = /* LUT   14 20  5 */ n866 ? n396 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n396 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2143 = /* LUT   17 20  2 */ n528 ? 1'b0 : 1'b1;
assign n1488 = /* LUT   19 18  3 */ n1370 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1430 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1430 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2145 = /* LUT   23 15  5 */ n158 ? 1'b1 : 1'b0;
assign n1665 = /* LUT   21 16  5 */ n1172 ? n1336 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1336 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n2147 = /* LUT   21 11  4 */ n35 ? 1'b1 : 1'b0;
assign n2148 = /* LUT   18 22  5 */ n272 ? io_0_25_1 ? n1259 ? n1025 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0;
assign n2149 = /* LUT   17  9  4 */ n1053 ? 1'b1 : 1'b0;
assign n2150 = /* LUT   11 19  1 */ n266 ? 1'b0 : 1'b1;
assign n2151 = /* LUT   10  9  1 */ n150 ? n195 ? n197 ? 1'b0 : n279 ? 1'b0 : 1'b1 : n197 ? n279 ? 1'b0 : 1'b1 : 1'b0 : n195 ? 1'b1 : 1'b0;
assign n2152 = /* LUT   22 15  1 */ n59 ? 1'b0 : n802 ? n244 ? n238 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2153 = /* LUT   13 17  7 */ n385 ? 1'b0 : n386 ? 1'b0 : n183 ? n256 ? 1'b0 : 1'b1 : 1'b0;
assign n2154 = /* LUT   18 21  1 */ n61 ? n1127 ? n899 ? 1'b1 : n731 ? 1'b1 : 1'b0 : n899 ? 1'b1 : 1'b0 : n1127 ? n899 ? n731 ? 1'b0 : 1'b1 : 1'b0 : n899 ? 1'b1 : 1'b0;
assign n2155 = /* LUT   19 14  6 */ n1319 ? n677 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n677 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2156 = /* LUT   16 13  2 */ n59 ? n244 ? 1'b0 : n440 ? n180 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2157 = /* LUT    5 18  0 */ n93 ? n52 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n52 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2158 = /* LUT   10 20  4 */ n140 ? 1'b1 : 1'b0;
assign n2159 = /* LUT   18  7  0 */ n1154 ? 1'b1 : 1'b0;
assign n1657 = /* LUT   21 15  1 */ n1574 ? n1543 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1543 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2161 = /* LUT   20 25  1 */ n212 ? 1'b1 : 1'b0;
assign n2162 = /* LUT   19 19  0 */ n159 ? 1'b1 : 1'b0;
assign n2163 = /* LUT   23 12  4 */ n35 ? 1'b1 : 1'b0;
assign n2164 = /* LUT   21 17  6 */ n1589 ? n1485 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1485 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2165 = /* LUT   21 12  5 */ n158 ? 1'b1 : 1'b0;
assign n2166 = /* LUT   18 25  4 */ n1417 ? n1387 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1387 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2167 = /* LUT   17 10  5 */ n32 ? 1'b1 : 1'b0;
assign n489  = /* LUT   11 16  0 */ n481 ? io_0_27_1 ? n355 ? 1'b0 : n340 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2169 = /* LUT   22 14  6 */ n140 ? 1'b1 : 1'b0;
assign n2170 = /* LUT   13 18  6 */ n185 ? 1'b0 : 1'b1;
assign n2171 = /* LUT   18 20  2 */ n1246 ? n1386 ? n709 ? 1'b1 : 1'b0 : n1247 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1386 ? 1'b0 : n1247 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n2172 = /* LUT   23 16  2 */ n44 ? 1'b1 : 1'b0;
assign n2173 = /* LUT   11 14  3 */ n453 ? n434 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n434 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n2174 = /* LUT   16  7  4 */ n1051 ? n904 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n904 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2175 = /* LUT   19 15  5 */ n212 ? 1'b1 : 1'b0;
assign n2176 = /* LUT   16 12  5 */ n770 ? 1'b0 : n159 ? 1'b1 : 1'b0;
assign n2177 = /* LUT   15 26  2 */ n1046 ? n882 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n882 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2178 = /* LUT   12 12  4 */ n36 ? 1'b1 : 1'b0;
assign n2179 = /* LUT   14 22  3 */ n158 ? 1'b1 : 1'b0;
assign n2180 = /* LUT   17 22  0 */ n979 ? 1'b0 : 1'b1;
assign n2182 = /* LUT   19 16  1 */ n212 ? 1'b1 : 1'b0;
assign n2183 = /* LUT   22 10  3 */ n1703 ? n1624 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n1624 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2184 = /* LUT    7 11  6 */ n66 ? n75 ? n80 ? 1'b1 : n107 ? 1'b1 : 1'b0 : n107 ? 1'b1 : 1'b0 : n75 ? n80 ? 1'b1 : 1'b0 : 1'b0;
assign n2185 = /* LUT   21 18  7 */ n1368 ? n1675 ? n575 ? 1'b1 : 1'b0 : n575 ? n812 ? 1'b1 : 1'b0 : 1'b1 : n1675 ? 1'b0 : n575 ? n812 ? 1'b1 : 1'b0 : 1'b1;
assign n2186 = /* LUT   21 13  6 */ n962 ? n1645 ? n575 ? 1'b1 : 1'b0 : n787 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1645 ? 1'b0 : n787 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2187 = /* LUT   12 15  6 */ n500 ? 1'b0 : 1'b1;
assign n2188 = /* LUT   18 24  7 */ n1278 ? n709 ? n930 ? 1'b0 : 1'b1 : n1276 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1276 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n907  = /* LUT   15  7  3 */ n904 ? 1'b0 : n900 ? n901 ? n903 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2189 = /* LUT   13 19  1 */ n268 ? 1'b0 : 1'b1;
assign n2190 = /* LUT   15 21  0 */ n1004 ? 1'b0 : 1'b1;
assign n2191 = /* LUT   18 23  3 */ n895 ? n1127 ? n55 ? 1'b1 : n731 ? 1'b0 : 1'b1 : 1'b1 : n1127 ? n55 ? n731 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2192 = /* LUT   23 17  5 */ n35 ? 1'b1 : 1'b0;
assign n2193 = /* LUT   11 15  0 */ n458 ? n303 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n303 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n2194 = /* LUT   19 12  4 */ n769 ? io_0_25_1 ? n59 ? 1'b0 : n802 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2195 = /* LUT    9 19  2 */ n257 ? n181 ? io_0_25_1 ? 1'b1 : 1'b0 : 1'b0 : n181 ? io_0_25_1 ? 1'b1 : 1'b0 : io_0_25_1 ? n258 ? 1'b0 : 1'b1 : 1'b0;
assign n2196 = /* LUT   12 19  5 */ n158 ? 1'b1 : 1'b0;
assign n2197 = /* LUT   14 17  2 */ n187 ? 1'b0 : n513 ? 1'b0 : n515 ? 1'b0 : n188 ? 1'b0 : 1'b1;
assign n2198 = /* LUT   17 12  6 */ n939 ? n1160 ? 1'b1 : n575 ? 1'b1 : 1'b0 : n1160 ? n575 ? 1'b0 : 1'b1 : 1'b0;
assign n2199 = /* LUT   17 23  7 */ n990 ? 1'b0 : 1'b1;
assign n2200 = /* LUT   22 21  1 */ n212 ? 1'b1 : 1'b0;
assign n1680 = /* LUT   21 19  0 */ n1610 ? n709 ? n930 ? 1'b0 : 1'b1 : n1471 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1471 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2204 = /* LUT   21 14  7 */ n1185 ? n1650 ? n575 ? 1'b1 : 1'b0 : n1547 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1650 ? 1'b0 : n1547 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2205 = /* LUT    9 16  4 */ io_0_20_0 ? 1'b0 : io_0_16_0 ? 1'b0 : io_25_0_0 ? 1'b0 : 1'b1;
assign n2206 = /* LUT   12 14  5 */ n473 ? 1'b0 : 1'b1;
assign n2207 = /* LUT   10 10  4 */ n290 ? n200 ? n150 ? 1'b0 : 1'b1 : n150 ? 1'b1 : 1'b0 : n200 ? 1'b1 : 1'b0;
assign n2208 = /* LUT   16 23  3 */ io_0_12_0 ? 1'b1 : 1'b0;
assign n2211 = /* LUT   13 20  0 */ n398 ? 1'b0 : 1'b1;
assign n2212 = /* LUT   15 10  1 */ n922 ? 1'b1 : 1'b0;
assign n2213 = /* LUT   20 19  2 */ n44 ? 1'b1 : 1'b0;
assign n2214 = /* LUT   11 12  1 */ n425 ? 1'b1 : 1'b0;
assign n2217 = /* LUT   19 13  3 */ n1305 ? n1444 ? n1437 ? n709 ? 1'b0 : 1'b1 : 1'b1 : n1437 ? 1'b0 : 1'b1 : n1444 ? n1437 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n1437 ? 1'b0 : n709 ? 1'b1 : 1'b0;
assign n2218 = /* LUT   16 10  7 */ n909 ? 1'b1 : 1'b0;
assign n2219 = /* LUT   15 24  0 */ n1026 ? n886 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n886 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2220 = /* LUT   12 18  6 */ n615 ? n500 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n500 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2221 = /* LUT   17 13  5 */ n784 ? n575 ? n1180 ? 1'b0 : 1'b1 : n951 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n951 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2222 = /* LUT   14 16  1 */ n699 ? 1'b1 : 1'b0;
assign n2223 = /* LUT   17 16  6 */ n1102 ? n1214 ? n709 ? 1'b1 : 1'b0 : n709 ? n1089 ? 1'b1 : 1'b0 : 1'b1 : n1214 ? 1'b0 : n709 ? n1089 ? 1'b1 : 1'b0 : 1'b1;
assign n1740 = /* LUT   22 20  2 */ n723 ? n721 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n721 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2225 = /* LUT   10 14  1 */ n213 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0;
assign n2226 = /* LUT   21 20  1 */ n212 ? 1'b1 : 1'b0;
assign n2229 = /* LUT    9 17  7 */ n42 ? 1'b1 : 1'b0;
assign n2230 = /* LUT   12 13  4 */ n35 ? 1'b1 : 1'b0;
assign n2231 = /* LUT   20 12  0 */ n159 ? 1'b1 : 1'b0;
assign n2232 = /* LUT   10 13  5 */ n310 ? n209 ? 1'b0 : n120 ? 1'b0 : 1'b1 : n209 ? n120 ? 1'b0 : 1'b1 : 1'b0;
assign n2233 = /* LUT   16 22  0 */ n1127 ? n891 ? n27 ? 1'b1 : n731 ? 1'b0 : 1'b1 : n27 ? n731 ? 1'b1 : 1'b0 : 1'b0 : n891 ? 1'b1 : 1'b0;
assign n2234 = /* LUT   10 16  5 */ n350 ? n235 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n235 ? 1'b1 : 1'b0;
assign n2235 = /* LUT   13 21  3 */ n183 ? 1'b0 : n179 ? n374 ? n495 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2236 = /* LUT   20 18  1 */ n159 ? 1'b1 : 1'b0;
assign n2237 = /* LUT   11 13  6 */ n159 ? 1'b1 : 1'b0;
assign n2238 = /* LUT   19 10  2 */ n44 ? 1'b1 : 1'b0;
assign n2239 = /* LUT   15 25  7 */ n1042 ? n897 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n897 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2240 = /* LUT    7 13  5 */ n122 ? n75 ? n80 ? 1'b0 : n124 ? 1'b1 : 1'b0 : 1'b0 : n75 ? n80 ? 1'b1 : n124 ? 1'b1 : 1'b0 : 1'b1;
assign n2241 = /* LUT   12 17  7 */ n603 ? n491 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n491 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2242 = /* LUT   14 19  0 */ n835 ? n269 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n269 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2243 = /* LUT   17 14  4 */ n1078 ? n1197 ? n575 ? 1'b1 : 1'b0 : n806 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1197 ? 1'b0 : n806 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n1221 = /* LUT   17 17  5 */ n984 ? 1'b0 : n1219 ? 1'b0 : 1'b1;
assign n2245 = /* LUT   22 23  3 */ n42 ? 1'b1 : 1'b0;
assign n2246 = /* LUT   21 21  2 */ n1611 ? n1696 ? n709 ? 1'b1 : 1'b0 : n1612 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1696 ? 1'b0 : n1612 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n407  = /* LUT   11  9  3 */ n195 ? n201 ? 1'b0 : n194 ? n200 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2247 = /* LUT   16 21  1 */ n42 ? 1'b1 : 1'b0;
assign n2248 = /* LUT   10 19  4 */ n35 ? 1'b1 : 1'b0;
assign n2249 = /* LUT   13 22  2 */ n400 ? 1'b0 : 1'b1;
assign n2250 = /* LUT    6 12  1 */ n68 ? 1'b1 : n70 ? 1'b1 : 1'b0;
assign n2251 = /* LUT   20 17  0 */ n1469 ? n1591 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1591 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2252 = /* LUT   23 20  6 */ n140 ? 1'b1 : 1'b0;
assign n2253 = /* LUT   11 10  7 */ n282 ? n154 ? n284 ? 1'b0 : 1'b1 : 1'b0 : n292 ? 1'b1 : 1'b0;
assign n2254 = /* LUT   19 11  1 */ n212 ? 1'b1 : 1'b0;
assign n2255 = /* LUT   12 16  0 */ n581 ? 1'b1 : 1'b0;
assign n1206 = /* LUT   17 15  3 */ n1204 ? n575 ? n1180 ? 1'b0 : 1'b1 : n976 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n976 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2257 = /* LUT   19 25  2 */ n44 ? 1'b1 : 1'b0;
assign n1715 = /* LUT   22 13  6 */ n1712 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1637 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1637 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2261 = /* LUT    7 15  2 */ n126 ? n84 ? 1'b0 : 1'b1 : n84 ? 1'b1 : 1'b0;
assign n2262 = /* LUT   21 22  3 */ n1411 ? n1699 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1699 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2263 = /* LUT   11 22  2 */ n44 ? 1'b1 : 1'b0;
assign n2264 = /* LUT   16 15  7 */ n769 ? n1099 ? io_0_25_1 ? n59 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2265 = /* LUT   10 15  7 */ n338 ? n226 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n226 ? 1'b1 : 1'b0;
assign n2266 = /* LUT   16 20  6 */ n781 ? n59 ? 1'b0 : 1'b1 : 1'b0;
assign n2267 = /* LUT   15 18  5 */ n158 ? 1'b1 : 1'b0;
assign n1324 = /* LUT   18 14  0 */ n1192 ? n705 ? n595 ? n1217 ? 1'b0 : 1'b1 : 1'b0 : n595 ? 1'b0 : 1'b1 : n705 ? n595 ? n1217 ? 1'b0 : 1'b1 : 1'b1 : n595 ? 1'b0 : 1'b1;
assign n2269 = /* LUT   20 16  7 */ n218 ? 1'b1 : 1'b0;
assign n2270 = /* LUT   12 20  5 */ n158 ? 1'b1 : 1'b0;
assign n2271 = /* LUT   11 11  4 */ n419 ? n280 ? 1'b0 : n282 ? 1'b0 : 1'b1 : n280 ? n282 ? 1'b0 : 1'b1 : 1'b0;
assign n1737 = /* LUT   22 18  1 */ n1671 ? n1736 ? n705 ? 1'b0 : 1'b1 : 1'b0 : n1662 ? 1'b1 : n705 ? 1'b1 : 1'b0;
assign n2273 = /* LUT   13  9  2 */ n552 ? 1'b1 : 1'b0;
assign n2274 = /* LUT   21 10  6 */ n1625 ? n1630 ? n1540 ? 1'b0 : n1538 ? 1'b0 : 1'b1 : n1538 ? 1'b0 : 1'b1 : n1630 ? n1540 ? 1'b0 : n1538 ? 1'b1 : 1'b0 : n1538 ? 1'b1 : 1'b0;
assign n2277 = /* LUT   17  8  2 */ n1156 ? 1'b1 : 1'b0;
assign n2278 = /* LUT   19 22  3 */ n1513 ? n1392 ? 1'b0 : n1258 ? 1'b0 : 1'b1 : n1392 ? n1258 ? 1'b0 : 1'b1 : 1'b0;
assign n2279 = /* LUT   22 17  5 */ n1638 ? n1732 ? n709 ? 1'b1 : 1'b0 : n1594 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1732 ? 1'b0 : n1594 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n2280 = /* LUT   16 16  3 */ n42 ? 1'b1 : 1'b0;
assign n2281 = /* LUT   22 12  5 */ n158 ? 1'b1 : 1'b0;
assign n946  = /* LUT   15 13  1 */ n779 ? n945 ? n689 ? n937 ? 1'b0 : 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2282 = /* LUT   20 20  4 */ n35 ? 1'b1 : 1'b0;
assign n2283 = /* LUT   16 14  4 */ n948 ? n937 ? 1'b0 : n244 ? 1'b0 : 1'b1 : 1'b0;
assign n2284 = /* LUT   16 19  7 */ n212 ? 1'b1 : 1'b0;
assign n2285 = /* LUT   15 19  6 */ n140 ? 1'b1 : 1'b0;
assign n2286 = /* LUT   15 14  5 */ n591 ? n770 ? 1'b0 : n163 ? n771 ? 1'b0 : 1'b1 : 1'b0 : n771 ? 1'b1 : 1'b0;
assign n1352 = /* LUT   18 17  1 */ n1216 ? n1227 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1227 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2288 = /* LUT   20 23  6 */ n42 ? 1'b1 : 1'b0;
assign n2289 = /* LUT   24 16  2 */ n218 ? 1'b1 : 1'b0;
assign n2290 = /* LUT   21 11  1 */ n212 ? 1'b1 : 1'b0;
assign n2293 = /* LUT   19 23  0 */ n1025 ? io_0_25_1 ? n272 ? n1024 ? 1'b1 : 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n1725 = /* LUT   22 16  6 */ n965 ? n1724 ? n575 ? 1'b1 : 1'b0 : n788 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1724 ? 1'b0 : n788 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2295 = /* LUT   22 15  4 */ n590 ? n802 ? n244 ? n59 ? 1'b0 : 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2296 = /* LUT   20 11  5 */ n140 ? 1'b1 : 1'b0;
assign n2297 = /* LUT   19 24  6 */ n1531 ? n796 ? 1'b0 : n1501 ? 1'b0 : 1'b1 : n796 ? n1501 ? 1'b0 : 1'b1 : 1'b0;
assign n2298 = /* LUT   11 20  0 */ n247 ? 1'b0 : 1'b1;
assign n2299 = /* LUT   16 13  5 */ n180 ? 1'b0 : n932 ? 1'b0 : n244 ? 1'b0 : n590 ? 1'b1 : 1'b0;
assign n2300 = /* LUT   16 18  4 */ n35 ? 1'b1 : 1'b0;
assign n2301 = /* LUT   10 20  1 */ n42 ? 1'b1 : 1'b0;
assign n2302 = /* LUT   15 16  7 */ n180 ? n972 ? n59 ? n244 ? 1'b0 : 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2303 = /* LUT   21 15  6 */ n1178 ? n1556 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1556 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2304 = /* LUT   15 15  6 */ n140 ? 1'b1 : 1'b0;
assign n2305 = /* LUT   18 16  2 */ n1343 ? n595 ? 1'b0 : n712 ? 1'b1 : 1'b0 : n595 ? n712 ? 1'b1 : 1'b0 : 1'b0;
assign n2306 = /* LUT    6  9  6 */ n66 ? 1'b0 : n107 ? 1'b1 : 1'b0;
assign n2307 = /* LUT   20 22  5 */ n1127 ? n1273 ? n697 ? n731 ? 1'b1 : 1'b0 : 1'b1 : n697 ? n731 ? 1'b0 : 1'b1 : 1'b0 : n1273 ? n697 ? 1'b0 : 1'b1 : n697 ? 1'b1 : 1'b0;
assign n2310 = /* LUT   24 15  3 */ n218 ? 1'b1 : 1'b0;
assign n675  = /* LUT   13 11  4 */ n557 ? n559 ? n569 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2311 = /* LUT   21 12  0 */ n159 ? 1'b1 : 1'b0;
assign n2312 = /* LUT   12 21  3 */ n520 ? 1'b0 : 1'b1;
assign n2313 = /* LUT   17 10  0 */ n712 ? n575 ? n930 ? 1'b0 : 1'b1 : n930 ? 1'b1 : 1'b0 : 1'b0;
assign n2314 = /* LUT   19 20  1 */ n272 ? n1377 ? io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0;
assign n2315 = /* LUT   22 19  7 */ n1734 ? n1693 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1693 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2316 = /* LUT   22 14  3 */ n42 ? 1'b1 : 1'b0;
assign n2317 = /* LUT   23 16  5 */ n158 ? 1'b1 : 1'b0;
assign n2318 = /* LUT   11 14  6 */ n456 ? n437 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n437 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n1070 = /* LUT   16 12  2 */ n778 ? n689 ? n943 ? 1'b0 : n779 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2320 = /* LUT   16 17  5 */ n158 ? 1'b1 : 1'b0;
assign n2321 = /* LUT   13 15  1 */ n577 ? 1'b1 : 1'b0;
assign n2322 = /* LUT   15 17  0 */ n159 ? 1'b1 : 1'b0;
assign n2323 = /* LUT   15 12  7 */ n125 ? 1'b1 : 1'b0;
assign n2324 = /* LUT   18 19  3 */ n1249 ? n820 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n820 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2325 = /* LUT   20 21  4 */ n1498 ? n1508 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1508 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2326 = /* LUT   24 14  0 */ n159 ? 1'b1 : 1'b0;
assign n2327 = /* LUT   13 12  5 */ n682 ? n569 ? 1'b0 : 1'b1 : n569 ? 1'b1 : 1'b0;
assign n2328 = /* LUT   21 13  3 */ n1554 ? n1644 ? n1438 ? n709 ? 1'b0 : 1'b1 : 1'b1 : n1438 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n1644 ? n1438 ? 1'b0 : 1'b1 : n1438 ? 1'b0 : n709 ? 1'b1 : 1'b0;
assign n2329 = /* LUT   19 21  6 */ n1025 ? 1'b0 : n641 ? n1502 ? 1'b1 : 1'b0 : n1398 ? 1'b1 : 1'b0;
assign n497  = /* LUT   11 17  4 */ n258 ? 1'b0 : n496 ? n374 ? 1'b0 : 1'b1 : 1'b1;
assign n2330 = /* LUT   24 17  6 */ n140 ? 1'b1 : 1'b0;
assign n2331 = /* LUT   15 21  5 */ n1001 ? 1'b0 : 1'b1;
assign n2332 = /* LUT   20  9  7 */ n1425 ? 1'b0 : n1294 ? 1'b1 : 1'b0;
assign n2333 = /* LUT   23 17  2 */ n1726 ? n1745 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1745 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2334 = /* LUT   11 15  5 */ n478 ? n300 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n300 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n2335 = /* LUT   11 18  6 */ n509 ? 1'b0 : 1'b1;
assign n2336 = /* LUT   16 11  3 */ n42 ? 1'b1 : 1'b0;
assign n2337 = /* LUT   13 16  0 */ n44 ? 1'b1 : 1'b0;
assign n2340 = /* LUT   18  9  5 */ n1283 ? 1'b1 : 1'b0;
assign n2341 = /* LUT   18 18  4 */ n1361 ? n1320 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1320 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2342 = /* LUT    6 11  4 */ n116 ? n71 ? 1'b0 : n81 ? 1'b0 : 1'b1 : n71 ? n81 ? 1'b0 : 1'b1 : 1'b0;
assign n2343 = /* LUT   14 10  0 */ n564 ? 1'b1 : 1'b0;
assign n2344 = /* LUT   19 17  3 */ n608 ? n709 ? n930 ? 1'b0 : 1'b1 : n1317 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1317 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2345 = /* LUT   22 21  4 */ n35 ? 1'b1 : 1'b0;
assign n2346 = /* LUT   24 13  1 */ n158 ? 1'b1 : 1'b0;
assign n2347 = /* LUT   13 13  6 */ n425 ? 1'b1 : 1'b0;
assign n2348 = /* LUT   21 14  2 */ n159 ? 1'b1 : 1'b0;
assign n2349 = /* LUT    9 16  3 */ io_25_0_0 ? 1'b0 : io_0_16_0 ? 1'b0 : io_0_20_0 ? 1'b0 : 1'b1;
assign n2350 = /* LUT   14 20  1 */ n862 ? n397 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n397 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2351 = /* LUT   19 18  7 */ n1174 ? n1338 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1338 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n2352 = /* LUT   10 10  1 */ n287 ? 1'b1 : 1'b0;
assign n2353 = /* LUT   16 23  6 */ n469 ? 1'b1 : 1'b0;
assign n1663 = /* LUT   21 16  1 */ n1646 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1290 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1290 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2355 = /* LUT   15 10  4 */ n918 ? 1'b1 : 1'b0;
assign n2356 = /* LUT   11 12  4 */ n424 ? 1'b1 : 1'b0;
assign n2357 = /* LUT   11 19  5 */ n262 ? 1'b0 : 1'b1;
assign n2358 = /* LUT   16 10  0 */ n914 ? 1'b1 : 1'b0;
assign n2359 = /* LUT    9 12  5 */ n203 ? 1'b0 : n204 ? 1'b1 : 1'b0;
assign n711  = /* LUT   13 17  3 */ n708 ? n710 ? n707 ? n706 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2360 = /* LUT   18 21  5 */ n888 ? n1127 ? n48 ? 1'b1 : n731 ? 1'b0 : 1'b1 : 1'b1 : n1127 ? n48 ? n731 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2361 = /* LUT   19 14  2 */ n1316 ? n1450 ? n575 ? 1'b1 : 1'b0 : n1448 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1450 ? 1'b0 : n1448 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2362 = /* LUT   22 20  7 */ n1486 ? n819 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n819 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2363 = /* LUT   16 24  4 */ io_4_33_1 ? 1'b1 : 1'b0;
assign n2364 = /* LUT    9 17  0 */ n141 ? n244 ? 1'b0 : n59 ? 1'b0 : n180 ? 1'b0 : 1'b1 : 1'b0;
assign n2365 = /* LUT   20 12  5 */ n158 ? 1'b1 : 1'b0;
assign n2366 = /* LUT   19 19  4 */ n158 ? 1'b1 : 1'b0;
assign n2367 = /* LUT   10 13  0 */ n305 ? n203 ? 1'b0 : n120 ? 1'b0 : 1'b1 : n203 ? n120 ? 1'b0 : 1'b1 : 1'b0;
assign n2368 = /* LUT   16 22  5 */ io_0_25_1 ? 1'b0 : 1'b1;
assign n2369 = /* LUT   22 11  0 */ n1708 ? n1627 ? 1'b0 : 1'b1 : n1627 ? 1'b1 : 1'b0;
assign n2370 = /* LUT   21 17  2 */ n1587 ? n1597 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1597 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2371 = /* LUT   20 15  1 */ n238 ? n180 ? 1'b0 : n932 ? 1'b0 : n244 ? 1'b0 : 1'b1 : 1'b0;
assign n2372 = /* LUT   11 13  3 */ n158 ? 1'b1 : 1'b0;
assign n2373 = /* LUT   11 16  4 */ n358 ? n83 ? n343 ? 1'b0 : 1'b1 : n343 ? n51 ? 1'b0 : 1'b1 : 1'b1 : n83 ? 1'b0 : n51 ? 1'b0 : 1'b1;
assign n2374 = /* LUT   16  9  1 */ n218 ? 1'b1 : 1'b0;
assign n2375 = /* LUT   13 18  2 */ n386 ? 1'b0 : 1'b1;
assign n2376 = /* LUT   15 20  3 */ n838 ? 1'b0 : 1'b1;
assign n2377 = /* LUT   18 20  6 */ n35 ? 1'b1 : 1'b0;
assign n2378 = /* LUT   16  7  0 */ n733 ? n900 ? 1'b0 : n737 ? 1'b0 : 1'b1 : n900 ? n737 ? 1'b0 : 1'b1 : 1'b0;
assign n1463 = /* LUT   19 15  1 */ n1461 ? n1459 ? 1'b1 : n1180 ? 1'b1 : 1'b0 : n1459 ? n1180 ? 1'b0 : 1'b1 : 1'b0;
assign n2381 = /* LUT   22 23  6 */ n140 ? 1'b1 : 1'b0;
assign n2382 = /* LUT   24 22  4 */ n1025 ? io_11_33_1 ? 1'b1 : 1'b0 : 1'b1;
assign n2383 = /* LUT    9 18  1 */ n158 ? 1'b1 : 1'b0;
assign n2384 = /* LUT   12 12  0 */ n429 ? 1'b1 : 1'b0;
assign n2385 = /* LUT   19 16  5 */ n158 ? 1'b1 : 1'b0;
assign n2386 = /* LUT   16 21  4 */ n140 ? 1'b1 : 1'b0;
assign n2387 = /* LUT   16 26  5 */ n44 ? 1'b1 : 1'b0;
assign n1674 = /* LUT   21 18  3 */ n1595 ? n575 ? n1180 ? 1'b0 : 1'b1 : n245 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n245 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2389 = /* LUT   15  7  7 */ n737 ? 1'b1 : n740 ? io_33_1_1 ? 1'b1 : 1'b0 : 1'b0;
assign n1413 = /* LUT   18 24  3 */ n1272 ? n1262 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1262 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2391 = /* LUT   20 14  2 */ n712 ? n1568 ? 1'b1 : 1'b0 : n1565 ? 1'b1 : 1'b0;
assign n2392 = /* LUT   23 20  1 */ n212 ? 1'b1 : 1'b0;
assign n413  = /* LUT   11 10  2 */ n280 ? 1'b0 : n296 ? 1'b0 : n281 ? 1'b0 : n295 ? 1'b0 : 1'b1;
assign n2394 = /* LUT    9 14  7 */ n156 ? n207 ? 1'b0 : n216 ? n206 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2395 = /* LUT   13 19  5 */ n515 ? 1'b0 : 1'b1;
assign n2396 = /* LUT   18 23  7 */ n897 ? n1127 ? n29 ? 1'b1 : n731 ? 1'b0 : 1'b1 : 1'b1 : n1127 ? n29 ? n731 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2397 = /* LUT   14 18  4 */ n831 ? n183 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n183 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2398 = /* LUT   14  7  3 */ n743 ? n649 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n649 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2399 = /* LUT   19 12  0 */ n948 ? n802 ? n59 ? 1'b0 : n244 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2400 = /* LUT   22 22  1 */ 1'b0 ? 1'b1 : 1'b0;
assign n2401 = /* LUT   12 19  1 */ n212 ? 1'b1 : 1'b0;
assign n2402 = /* LUT   17 12  2 */ n1063 ? n1182 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1182 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2403 = /* LUT   10 15  2 */ n333 ? n221 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n221 ? 1'b1 : 1'b0;
assign n2404 = /* LUT   16 20  3 */ n238 ? n244 ? 1'b0 : n937 ? 1'b0 : 1'b1 : 1'b0;
assign n1683 = /* LUT   21 19  4 */ n1562 ? n1682 ? n709 ? 1'b1 : 1'b0 : n1592 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1682 ? 1'b0 : n1592 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n2408 = /* LUT   15  9  1 */ n917 ? 1'b1 : 1'b0;
assign n2409 = /* LUT   18 14  5 */ n1093 ? n1326 ? n709 ? n1067 ? 1'b1 : 1'b0 : 1'b0 : 1'b1 : n1326 ? n709 ? n1067 ? 1'b1 : 1'b0 : 1'b0 : n709 ? 1'b0 : 1'b1;
assign n1558 = /* LUT   20 13  3 */ n1441 ? n1542 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1542 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2411 = /* LUT   11 11  1 */ n416 ? n283 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n283 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2412 = /* LUT   22 18  6 */ n1245 ? n1739 ? n595 ? 1'b0 : n705 ? 1'b0 : 1'b1 : n595 ? 1'b0 : 1'b1 : n1739 ? n595 ? n705 ? 1'b1 : 1'b0 : n705 ? 1'b0 : 1'b1 : n595 ? n705 ? 1'b1 : 1'b0 : 1'b1;
assign n2413 = /* LUT   10 17  2 */ n361 ? n241 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n241 ? 1'b1 : 1'b0;
assign n2414 = /* LUT    9 15  0 */ n162 ? n167 ? n164 ? n166 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2415 = /* LUT   13 20  4 */ n189 ? 1'b0 : 1'b1;
assign n2416 = /* LUT   18 13  1 */ n712 ? n1312 ? 1'b1 : 1'b0 : n953 ? 1'b1 : 1'b0;
assign n2417 = /* LUT   14 13  5 */ n158 ? 1'b1 : 1'b0;
assign n2418 = /* LUT   19 22  6 */ n1516 ? n1395 ? 1'b0 : n1258 ? 1'b0 : 1'b1 : n1395 ? n1258 ? 1'b0 : 1'b1 : 1'b0;
assign n2421 = /* LUT   19 13  7 */ n1171 ? n1321 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1321 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n1730 = /* LUT   22 17  0 */ n1669 ? n705 ? 1'b0 : n1668 ? 1'b1 : 1'b0 : n705 ? 1'b1 : n1582 ? 1'b1 : 1'b0;
assign n2423 = /* LUT   15 13  6 */ n770 ? 1'b0 : n35 ? 1'b1 : 1'b0;
assign n2424 = /* LUT   12 18  2 */ n611 ? n486 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n486 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2425 = /* LUT   14 16  5 */ n322 ? n807 ? 1'b1 : io_0_25_1 ? io_33_1_1 ? 1'b1 : 1'b0 : 1'b1 : n807 ? 1'b1 : io_0_25_1 ? io_33_1_1 ? 1'b1 : 1'b0 : 1'b0;
assign n1187 = /* LUT   17 13  1 */ n783 ? n575 ? n1180 ? 1'b0 : 1'b1 : n954 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n954 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2427 = /* LUT   16 19  2 */ n35 ? 1'b1 : 1'b0;
assign n2428 = /* LUT   21 20  5 */ n158 ? 1'b1 : 1'b0;
assign n955  = /* LUT   15 14  0 */ n782 ? n776 ? 1'b0 : n244 ? n591 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n1353 = /* LUT   18 17  4 */ n722 ? n1114 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1114 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2432 = /* LUT   18 26  5 */ n1421 ? n1282 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1282 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2433 = /* LUT   10 16  1 */ n346 ? n231 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n231 ? 1'b1 : 1'b0;
assign n2434 = /* LUT   13 21  7 */ n258 ? io_0_25_1 ? n181 ? 1'b0 : 1'b1 : 1'b1 : io_0_25_1 ? n257 ? n181 ? 1'b0 : 1'b1 : 1'b0 : 1'b1;
assign n2435 = /* LUT   18 12  2 */ n44 ? 1'b1 : 1'b0;
assign n2436 = /* LUT   14 12  6 */ n770 ? n774 ? n159 ? 1'b1 : 1'b0 : n28 ? 1'b1 : 1'b0 : n774 ? 1'b0 : n28 ? 1'b1 : 1'b0;
assign n2437 = /* LUT   19 23  5 */ n272 ? n1403 ? io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0;
assign n2438 = /* LUT   19 10  6 */ n140 ? 1'b1 : 1'b0;
assign n1723 = /* LUT   22 16  3 */ n1173 ? n1337 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1337 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n2440 = /* LUT   12 17  3 */ n599 ? n471 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n471 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2441 = /* LUT   14 19  4 */ n848 ? n187 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n187 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n1196 = /* LUT   17 14  0 */ n1080 ? n575 ? n1180 ? 1'b0 : 1'b1 : n975 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n975 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2443 = /* LUT   19 24  1 */ n1526 ? n1406 ? 1'b0 : n1501 ? 1'b0 : 1'b1 : n1406 ? n1501 ? 1'b0 : 1'b1 : 1'b0;
assign n2444 = /* LUT   16 18  1 */ n212 ? 1'b1 : 1'b0;
assign n2445 = /* LUT   21 21  6 */ n212 ? 1'b1 : 1'b0;
assign n2446 = /* LUT   13 25  0 */ n732 ? 1'b0 : n354 ? n374 ? 1'b0 : 1'b1 : 1'b1;
assign n2447 = /* LUT   15 15  3 */ n42 ? 1'b1 : 1'b0;
assign n2448 = /* LUT   10 19  0 */ n159 ? 1'b1 : 1'b0;
assign n2449 = /* LUT   13 11  1 */ n569 ? io_33_1_1 ? 1'b0 : 1'b1 : n674 ? n559 ? 1'b0 : io_33_1_1 ? 1'b0 : 1'b1 : io_33_1_1 ? 1'b0 : 1'b1;
assign n2450 = /* LUT   13 22  6 */ n401 ? 1'b0 : 1'b1;
assign n2451 = /* LUT   18 15  3 */ n814 ? n1333 ? n575 ? 1'b1 : 1'b0 : n483 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1333 ? 1'b0 : n483 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2452 = /* LUT   14 15  7 */ n358 ? n703 ? n771 ? 1'b1 : n770 ? 1'b1 : 1'b0 : n771 ? 1'b1 : 1'b0 : 1'b0;
assign n2453 = /* LUT   19 20  4 */ n1025 ? io_0_25_1 ? n1380 ? 1'b1 : n272 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2454 = /* LUT   19 11  5 */ n158 ? 1'b1 : 1'b0;
assign n2455 = /* LUT   22 19  2 */ n1676 ? n575 ? n1606 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n1606 ? 1'b1 : 1'b0 : 1'b0;
assign n2456 = /* LUT   17 15  7 */ n139 ? n575 ? n1180 ? 1'b0 : 1'b1 : n974 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n974 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2457 = /* LUT   16 17  0 */ n159 ? 1'b1 : 1'b0;
assign n2458 = /* LUT   22 13  2 */ n42 ? 1'b1 : 1'b0;
assign n2459 = /* LUT   15 12  2 */ n753 ? n762 ? 1'b1 : n152 ? 1'b1 : 1'b0 : n762 ? n152 ? 1'b0 : 1'b1 : 1'b0;
assign n2460 = /* LUT   18 19  6 */ n1375 ? n1229 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1229 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n1098 = /* LUT   16 15  3 */ n780 ? n943 ? n778 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2461 = /* LUT   23 13  5 */ n140 ? 1'b1 : 1'b0;
assign n2462 = /* LUT   24 14  5 */ n158 ? 1'b1 : 1'b0;
assign n2463 = /* LUT    9 10  3 */ io_4_0_0 ? n136 ? n75 ? 1'b0 : 1'b1 : 1'b1 : 1'b0;
assign n2467 = /* LUT   15 18  1 */ n212 ? 1'b1 : 1'b0;
assign n2468 = /* LUT   14 14  0 */ n770 ? 1'b0 : n218 ? 1'b1 : 1'b0;
assign n2469 = /* LUT   17 11  4 */ n1060 ? n1169 ? n709 ? 1'b0 : n930 ? 1'b0 : 1'b1 : n930 ? 1'b0 : 1'b1 : n1169 ? n709 ? n930 ? 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n709 ? 1'b1 : n930 ? 1'b0 : 1'b1;
assign n2470 = /* LUT   19 21  3 */ n641 ? n1146 ? n1025 ? 1'b0 : 1'b1 : 1'b0 : n1382 ? n1025 ? 1'b0 : 1'b1 : 1'b0;
assign n2471 = /* LUT   23 14  1 */ n212 ? 1'b1 : 1'b0;
assign n2472 = /* LUT   24 17  1 */ n212 ? 1'b1 : 1'b0;
assign n2473 = /* LUT   21 10  2 */ n1535 ? 1'b0 ? n1425 ? 1'b1 : 1'b0 : n1425 ? 1'b0 : 1'b1 : 1'b0 ? n1425 ? 1'b0 : 1'b1 : n1425 ? 1'b1 : 1'b0;
assign n2476 = /* LUT   22 12  1 */ n212 ? 1'b1 : 1'b0;
assign n2477 = /* LUT   13 16  7 */ n212 ? 1'b1 : 1'b0;
assign n2478 = /* LUT    7 12  7 */ n111 ? 1'b1 : n137 ? 1'b1 : n109 ? 1'b0 : n108 ? 1'b1 : 1'b0;
assign n1363 = /* LUT   18 18  1 */ n1224 ? n575 ? n1362 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n1362 ? 1'b1 : 1'b0 : 1'b0;
assign n2480 = /* LUT   20 20  0 */ n159 ? 1'b1 : 1'b0;
assign n2481 = /* LUT   23 18  3 */ n35 ? 1'b1 : 1'b0;
assign n2482 = /* LUT   14 10  5 */ n758 ? 1'b1 : 1'b0;
assign n2483 = /* LUT   16 14  0 */ n778 ? 1'b0 : n935 ? n943 ? n780 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2484 = /* LUT    5 17  6 */ n91 ? n50 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n50 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2485 = /* LUT   13 13  3 */ n431 ? 1'b0 : 1'b1;
assign n2486 = /* LUT   17 20  5 */ n396 ? 1'b0 : 1'b1;
assign n2487 = /* LUT   19 18  2 */ n1355 ? n1487 ? n575 ? 1'b1 : 1'b0 : n1468 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1487 ? 1'b0 : n1468 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2488 = /* LUT   23 15  2 */ n44 ? 1'b1 : 1'b0;
assign n2489 = /* LUT   21 16  4 */ n964 ? n1664 ? n575 ? 1'b1 : 1'b0 : n785 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1664 ? 1'b0 : n785 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2490 = /* LUT   21 11  5 */ n158 ? 1'b1 : 1'b0;
assign n2491 = /* LUT   18 22  6 */ n1025 ? n1260 ? io_0_25_1 ? 1'b1 : 1'b0 : io_0_25_1 ? n272 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2494 = /* LUT   10  9  0 */ n277 ? n150 ? n194 ? 1'b0 : n279 ? 1'b0 : 1'b1 : n194 ? 1'b1 : 1'b0 : n150 ? n194 ? n279 ? 1'b0 : 1'b1 : 1'b0 : n194 ? 1'b1 : 1'b0;
assign n2495 = /* LUT   22 15  0 */ n590 ? n244 ? 1'b0 : n525 ? 1'b0 : n59 ? 1'b1 : 1'b0 : 1'b0;
assign n2496 = /* LUT   13 17  4 */ n594 ? n711 ? n593 ? 1'b0 : io_0_25_1 ? 1'b1 : 1'b0 : io_0_25_1 ? 1'b1 : 1'b0 : io_0_25_1 ? 1'b1 : 1'b0;
assign n2497 = /* LUT   18 21  0 */ n731 ? n1127 ? n60 ? 1'b1 : 1'b0 : n898 ? 1'b1 : 1'b0 : n898 ? 1'b1 : 1'b0;
assign n2498 = /* LUT   20 11  1 */ n44 ? 1'b1 : 1'b0;
assign n2499 = /* LUT   16 13  1 */ n770 ? 1'b0 : n44 ? 1'b1 : 1'b0;
assign n2500 = /* LUT    5 18  7 */ n100 ? n29 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n29 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2501 = /* LUT   10 20  5 */ n218 ? 1'b1 : 1'b0;
assign n2502 = /* LUT   15 16  3 */ n59 ? n777 ? 1'b0 : n781 ? 1'b1 : 1'b0 : 1'b0;
assign n2503 = /* LUT   21 15  2 */ n1571 ? n1657 ? n930 ? 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? 1'b0 : 1'b1 : n1657 ? n930 ? n709 ? 1'b1 : 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? n709 ? 1'b1 : 1'b0 : 1'b1;
assign n2504 = /* LUT   20 25  0 */ n159 ? 1'b1 : 1'b0;
assign n2505 = /* LUT   17 21  6 */ n1243 ? n1240 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1240 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2506 = /* LUT   19 19  1 */ n44 ? 1'b1 : 1'b0;
assign n2509 = /* LUT   23 12  3 */ n42 ? 1'b1 : 1'b0;
assign n2510 = /* LUT   21 17  7 */ n140 ? 1'b1 : 1'b0;
assign n2511 = /* LUT   21 12  4 */ n35 ? 1'b1 : 1'b0;
assign n2512 = /* LUT   12 21  7 */ n523 ? 1'b0 : 1'b1;
assign n2513 = /* LUT   17 10  4 */ n32 ? 1'b1 : 1'b0;
assign n2514 = /* LUT   22 14  7 */ n218 ? 1'b1 : 1'b0;
assign n2515 = /* LUT   13 18  5 */ n345 ? 1'b0 : 1'b1;
assign n2516 = /* LUT   23 16  1 */ n212 ? 1'b1 : 1'b0;
assign n2517 = /* LUT   11 14  2 */ n452 ? n433 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n433 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n1072 = /* LUT   16 12  6 */ n59 ? 1'b1 : n440 ? 1'b0 : 1'b1;
assign n2518 = /* LUT    5 19  0 */ n101 ? n60 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n60 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2519 = /* LUT   22 24  0 */ n42 ? 1'b1 : 1'b0;
assign n2520 = /* LUT   15 17  4 */ n35 ? 1'b1 : 1'b0;
assign n2521 = /* LUT   20 24  7 */ n1409 ? n1621 ? n1620 ? n1410 ? 1'b1 : 1'b0 : 1'b0 : n1620 ? n1410 ? 1'b0 : 1'b1 : 1'b0 : n1621 ? n1620 ? 1'b0 : n1410 ? 1'b1 : 1'b0 : n1620 ? 1'b0 : n1410 ? 1'b0 : 1'b1;
assign n2522 = /* LUT   17 22  7 */ n983 ? 1'b0 : 1'b1;
assign n2523 = /* LUT   14 11  3 */ n659 ? 1'b1 : 1'b0;
assign n2524 = /* LUT   19 16  0 */ n159 ? 1'b1 : 1'b0;
assign n2525 = /* LUT   22 10  4 */ n1704 ? n1294 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n1294 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n1675 = /* LUT   21 18  6 */ n575 ? n1180 ? 1'b0 : 1'b1 : n1602 ? n825 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n825 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2527 = /* LUT   21 13  7 */ n1642 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1163 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1163 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2528 = /* LUT   12 15  1 */ n485 ? 1'b0 : 1'b1;
assign n2529 = /* LUT   15  7  0 */ n736 ? n902 ? n905 ? io_33_1_1 ? 1'b0 : 1'b1 : 1'b0 : io_33_1_1 ? 1'b0 : 1'b1 : io_33_1_1 ? 1'b0 : 1'b1;
assign n1414 = /* LUT   18 24  4 */ n1270 ? n1413 ? n709 ? n930 ? 1'b0 : 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n1413 ? n709 ? n930 ? 1'b0 : 1'b1 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2531 = /* LUT   13 19  2 */ n516 ? 1'b0 : 1'b1;
assign n2532 = /* LUT   15 21  1 */ n1005 ? 1'b0 : 1'b1;
assign n2533 = /* LUT   18 23  2 */ n731 ? n1127 ? n54 ? 1'b1 : 1'b0 : n894 ? 1'b1 : 1'b0 : n894 ? 1'b1 : 1'b0;
assign n1747 = /* LUT   23 17  6 */ n1721 ? n1718 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1718 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n2535 = /* LUT   11 15  1 */ n474 ? n304 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n304 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n2536 = /* LUT   16 11  7 */ n218 ? 1'b1 : 1'b0;
assign n2537 = /* LUT    5 20  1 */ io_0_28_1 ? 1'b0 : io_0_25_1 ? 1'b1 : 1'b0;
assign n2540 = /* LUT   18  9  1 */ n755 ? 1'b1 : 1'b0;
assign n2541 = /* LUT   12 19  4 */ n35 ? 1'b1 : 1'b0;
assign n2542 = /* LUT   17 23  0 */ n991 ? 1'b0 : 1'b1;
assign n2543 = /* LUT   22 21  0 */ n159 ? 1'b1 : 1'b0;
assign n1681 = /* LUT   21 19  1 */ n1069 ? n1680 ? n709 ? 1'b1 : 1'b0 : n1481 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1680 ? 1'b0 : n1481 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n1650 = /* LUT   21 14  6 */ n1577 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1180 ? n1634 ? 1'b0 : 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1180 ? n1634 ? 1'b0 : 1'b1 : 1'b1;
assign n2548 = /* LUT    9 16  7 */ n212 ? n218 ? n42 ? n158 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2549 = /* LUT   12 14  2 */ n470 ? 1'b0 : 1'b1;
assign n2552 = /* LUT   16 23  2 */ io_3_33_1 ? 1'b1 : 1'b0;
assign n2553 = /* LUT   13 20  3 */ n527 ? 1'b0 : 1'b1;
assign n2554 = /* LUT   15 10  0 */ n754 ? 1'b1 : 1'b0;
assign n2555 = /* LUT   20 19  5 */ n158 ? 1'b1 : 1'b0;
assign n2556 = /* LUT   11 12  0 */ n426 ? 1'b1 : 1'b0;
assign n2559 = /* LUT   16 10  4 */ n1056 ? 1'b1 : 1'b0;
assign n2560 = /* LUT    9 12  1 */ n155 ? n108 ? 1'b1 : n121 ? 1'b1 : n154 ? 1'b1 : 1'b0 : n108 ? 1'b0 : n121 ? 1'b0 : n154 ? 1'b1 : 1'b0;
assign n2561 = /* LUT   15 24  7 */ n1033 ? n891 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n891 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2562 = /* LUT   12 18  7 */ n616 ? n501 ? 1'b0 : 1'b1 : n501 ? 1'b1 : 1'b0;
assign n2563 = /* LUT   17 16  1 */ n977 ? n978 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n978 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n1741 = /* LUT   22 20  3 */ n1687 ? n1740 ? n930 ? 1'b0 : n709 ? 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n1740 ? n930 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n930 ? n709 ? 1'b0 : 1'b1 : 1'b1;
assign n2565 = /* LUT   10 14  2 */ n214 ? io_0_25_1 ? n213 ? 1'b0 : 1'b1 : 1'b1 : io_0_25_1 ? n213 ? 1'b1 : 1'b0 : 1'b0;
assign n2566 = /* LUT   16 24  0 */ io_7_33_0 ? 1'b1 : 1'b0;
assign n2567 = /* LUT   21 20  0 */ n159 ? 1'b1 : 1'b0;
assign n2570 = /* LUT   12 13  3 */ n42 ? 1'b1 : 1'b0;
assign n2571 = /* LUT   20 12  1 */ n212 ? 1'b1 : 1'b0;
assign n2572 = /* LUT   10 13  4 */ n309 ? n204 ? 1'b0 : n120 ? 1'b0 : 1'b1 : n204 ? n120 ? 1'b0 : 1'b1 : 1'b0;
assign n2573 = /* LUT   16 22  1 */ n731 ? n52 ? n1127 ? 1'b1 : n893 ? 1'b1 : 1'b0 : n1127 ? 1'b0 : n893 ? 1'b1 : 1'b0 : n893 ? 1'b1 : 1'b0;
assign n2574 = /* LUT   13 21  0 */ n719 ? n542 ? 1'b0 : 1'b1 : 1'b1;
assign n2575 = /* LUT   20 18  6 */ n44 ? 1'b1 : 1'b0;
assign n2576 = /* LUT   20 15  5 */ n238 ? n1578 ? n244 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2577 = /* LUT   11 13  7 */ n212 ? 1'b1 : 1'b0;
assign n655  = /* LUT   13  7  1 */ n648 ? n654 ? 1'b1 : 1'b0 : n652 ? 1'b1 : 1'b0;
assign n2579 = /* LUT   15 25  0 */ n1034 ? n893 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n893 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2580 = /* LUT   15 20  7 */ n842 ? 1'b0 : 1'b1;
assign n2581 = /* LUT   18 11  3 */ n218 ? 1'b1 : 1'b0;
assign n2582 = /* LUT   12 17  6 */ n602 ? n490 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n490 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2583 = /* LUT   17 17  2 */ n1107 ? n1220 ? n930 ? 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? 1'b0 : 1'b1 : n1220 ? n930 ? n709 ? 1'b1 : 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? n709 ? 1'b1 : 1'b0 : 1'b1;
assign n2584 = /* LUT   22 23  2 */ n44 ? 1'b1 : 1'b0;
assign n2585 = /* LUT   11  9  4 */ n65 ? 1'b0 : n407 ? n152 ? n151 ? 1'b0 : 1'b1 : 1'b1 : 1'b1;
assign n2586 = /* LUT   16 21  0 */ n44 ? 1'b1 : 1'b0;
assign n2587 = /* LUT   13 22  1 */ n399 ? 1'b0 : 1'b1;
assign n2588 = /* LUT   20 17  7 */ n42 ? 1'b1 : 1'b0;
assign n2589 = /* LUT   20 14  6 */ n1551 ? n709 ? n930 ? 1'b0 : 1'b1 : n1328 ? 1'b0 : n930 ? 1'b0 : 1'b1 : n709 ? n930 ? 1'b0 : 1'b1 : n1328 ? n930 ? 1'b1 : 1'b0 : 1'b1;
assign n2590 = /* LUT   23 20  5 */ n158 ? 1'b1 : 1'b0;
assign n2591 = /* LUT   14 18  0 */ n827 ? n385 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n385 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2594 = /* LUT   21 22  2 */ n1238 ? n1603 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1603 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2595 = /* LUT   11 22  5 */ n158 ? 1'b1 : 1'b0;
assign n1099 = /* LUT   16 15  6 */ n440 ? 1'b0 : n180 ? 1'b1 : 1'b0;
assign n2596 = /* LUT   10 15  6 */ n337 ? n225 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n225 ? 1'b1 : 1'b0;
assign n2597 = /* LUT   16 20  7 */ n238 ? n244 ? n525 ? 1'b0 : n59 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2598 = /* LUT   21 24  1 */ n158 ? 1'b1 : 1'b0;
assign n2599 = /* LUT   15 18  4 */ n35 ? 1'b1 : 1'b0;
assign n2600 = /* LUT   18 14  1 */ n1191 ? n1324 ? n705 ? 1'b0 : 1'b1 : n1202 ? 1'b1 : n705 ? 1'b1 : 1'b0 : n1324 ? 1'b0 : n1202 ? 1'b1 : n705 ? 1'b1 : 1'b0;
assign n2601 = /* LUT   20 16  0 */ n159 ? 1'b1 : 1'b0;
assign n2602 = /* LUT   12 20  6 */ n140 ? 1'b1 : 1'b0;
assign n2603 = /* LUT   20 13  7 */ n44 ? 1'b1 : 1'b0;
assign n2604 = /* LUT   11 11  5 */ n420 ? n281 ? 1'b0 : n282 ? 1'b0 : 1'b1 : n281 ? n282 ? 1'b0 : 1'b1 : 1'b0;
assign n2605 = /* LUT   22 18  2 */ n712 ? n1737 ? 1'b1 : 1'b0 : n1491 ? 1'b1 : 1'b0;
assign n2606 = /* LUT    9 15  4 */ n220 ? n223 ? n221 ? n222 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n1630 = /* LUT   21 10  5 */ n1425 ? n1629 ? n1623 ? n1536 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2609 = /* LUT   14 13  1 */ n212 ? 1'b1 : 1'b0;
assign n2610 = /* LUT   19 22  2 */ n1512 ? n1391 ? 1'b0 : n1258 ? 1'b0 : 1'b1 : n1391 ? n1258 ? 1'b0 : 1'b1 : 1'b0;
assign n1732 = /* LUT   22 17  4 */ n1727 ? n709 ? n930 ? 1'b0 : 1'b1 : n1660 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1660 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2612 = /* LUT   16 16  4 */ n35 ? 1'b1 : 1'b0;
assign n2613 = /* LUT    7 12  2 */ n78 ? 1'b0 : n77 ? 1'b0 : n79 ? 1'b1 : 1'b0;
assign n2614 = /* LUT   15 13  2 */ n782 ? n946 ? n777 ? n591 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2615 = /* LUT   20 20  5 */ n158 ? 1'b1 : 1'b0;
assign n1086 = /* LUT   16 14  5 */ n780 ? n778 ? n943 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2616 = /* LUT   16 19  6 */ n159 ? 1'b1 : 1'b0;
assign n2617 = /* LUT   15 19  7 */ n218 ? 1'b1 : 1'b0;
assign n2618 = /* LUT   18 17  0 */ n1115 ? n575 ? n824 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n824 ? 1'b1 : 1'b0 : 1'b0;
assign n2619 = /* LUT   15 14  4 */ n771 ? n770 ? n591 ? 1'b0 : 1'b1 : n591 ? 1'b1 : 1'b0 : n770 ? n591 ? 1'b0 : 1'b1 : 1'b0;
assign n2620 = /* LUT   19  9  0 */ n218 ? 1'b1 : 1'b0;
assign n2621 = /* LUT   21 11  2 */ n44 ? 1'b1 : 1'b0;
assign n2622 = /* LUT   18 12  6 */ n140 ? 1'b1 : 1'b0;
assign n2625 = /* LUT   14 12  2 */ n549 ? n764 ? 1'b1 : n152 ? 1'b0 : 1'b1 : n764 ? n152 ? 1'b1 : 1'b0 : 1'b0;
assign n2626 = /* LUT   19 23  1 */ n272 ? n1400 ? io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0;
assign n2627 = /* LUT   22 16  7 */ n1661 ? n1725 ? n1573 ? n709 ? 1'b0 : 1'b1 : 1'b1 : n1573 ? 1'b0 : 1'b1 : n1725 ? n1573 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n1573 ? 1'b0 : n709 ? 1'b1 : 1'b0;
assign n2628 = /* LUT   20 11  4 */ n158 ? 1'b1 : 1'b0;
assign n2629 = /* LUT   19 24  5 */ n1530 ? n1410 ? 1'b0 : n1501 ? 1'b0 : 1'b1 : n1410 ? n1501 ? 1'b0 : 1'b1 : 1'b0;
assign n2630 = /* LUT   11 20  7 */ n254 ? 1'b0 : 1'b1;
assign n2631 = /* LUT   16 13  4 */ n59 ? n244 ? 1'b0 : n440 ? n180 ? 1'b0 : 1'b1 : 1'b0 : n244 ? 1'b0 : n440 ? 1'b0 : n180 ? 1'b1 : 1'b0;
assign n2632 = /* LUT   16 18  5 */ n158 ? 1'b1 : 1'b0;
assign n972  = /* LUT   15 16  6 */ n540 ? n59 ? n440 ? 1'b0 : 1'b1 : n440 ? 1'b1 : 1'b0 : 1'b0;
assign n2633 = /* LUT   21 15  7 */ n35 ? 1'b1 : 1'b0;
assign n2634 = /* LUT   15 15  7 */ n218 ? 1'b1 : 1'b0;
assign n2635 = /* LUT   18 16  3 */ n1344 ? n705 ? 1'b0 : n712 ? 1'b1 : 1'b0 : n705 ? n712 ? 1'b1 : 1'b0 : 1'b0;
assign n2636 = /* LUT   20 22  2 */ n1025 ? n1504 ? 1'b1 : 1'b0 : n1618 ? n641 ? n1504 ? 1'b1 : 1'b0 : 1'b0 : n641 ? 1'b1 : 1'b0;
assign n2639 = /* LUT   24 15  2 */ n35 ? 1'b1 : 1'b0;
assign n2640 = /* LUT   13 11  5 */ n558 ? n675 ? n562 ? 1'b0 : io_33_1_1 ? 1'b1 : 1'b0 : n562 ? 1'b0 : 1'b1 : n675 ? n562 ? io_33_1_1 ? 1'b1 : 1'b0 : 1'b0 : n562 ? 1'b1 : 1'b0;
assign n2641 = /* LUT   21 12  3 */ n42 ? 1'b1 : 1'b0;
assign n2642 = /* LUT   12 21  2 */ n519 ? 1'b0 : 1'b1;
assign n2643 = /* LUT   19 20  0 */ n1025 ? io_0_25_1 ? n1376 ? 1'b1 : n272 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2644 = /* LUT   22 19  6 */ n1733 ? n1689 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1689 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2645 = /* LUT   23 16  4 */ n35 ? 1'b1 : 1'b0;
assign n2646 = /* LUT   11 21  0 */ n529 ? 1'b1 : 1'b0;
assign n1071 = /* LUT   16 12  3 */ n244 ? 1'b0 : n1070 ? n525 ? 1'b0 : n59 ? 1'b0 : 1'b1 : 1'b0;
assign n2648 = /* LUT   16 17  4 */ n35 ? 1'b1 : 1'b0;
assign n2649 = /* LUT   13 15  2 */ n696 ? 1'b1 : 1'b0;
assign n2650 = /* LUT   15 17  1 */ n212 ? 1'b1 : 1'b0;
assign n2651 = /* LUT   18 19  2 */ n1371 ? n815 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n815 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2652 = /* LUT   20 21  3 */ n35 ? 1'b1 : 1'b0;
assign n2653 = /* LUT   17 25  3 */ n1044 ? n1150 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1150 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2654 = /* LUT   23 13  1 */ n35 ? 1'b1 : 1'b0;
assign n2655 = /* LUT   24 14  1 */ n212 ? 1'b1 : 1'b0;
assign n2656 = /* LUT   13 12  4 */ n681 ? n568 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n568 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2657 = /* LUT   21 13  0 */ n1555 ? n575 ? n1553 ? 1'b1 : 1'b0 : 1'b0 : n575 ? n1458 ? 1'b1 : 1'b0 : 1'b1;
assign n2658 = /* LUT   17 11  0 */ n1167 ? n926 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n926 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2659 = /* LUT   19 21  7 */ n641 ? n1494 ? 1'b1 : n1025 ? 1'b1 : 1'b0 : n1397 ? 1'b1 : n1025 ? 1'b1 : 1'b0;
assign n2660 = /* LUT   11 17  5 */ n482 ? n497 ? n493 ? n344 ? 1'b1 : 1'b0 : 1'b0 : n493 ? 1'b1 : 1'b0 : 1'b0;
assign n2661 = /* LUT   23 14  5 */ n158 ? 1'b1 : 1'b0;
assign n2662 = /* LUT   24 17  5 */ n158 ? 1'b1 : 1'b0;
assign n2663 = /* LUT   15 21  6 */ n1002 ? 1'b0 : 1'b1;
assign n556  = /* LUT   12 10  2 */ n151 ? n410 ? 1'b1 : 1'b0 : n555 ? 1'b1 : 1'b0;
assign n1746 = /* LUT   23 17  3 */ n1720 ? n1717 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1717 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n2666 = /* LUT   11 18  1 */ n504 ? 1'b0 : 1'b1;
assign n2667 = /* LUT   16 11  2 */ n44 ? 1'b1 : 1'b0;
assign n2668 = /* LUT   13 16  3 */ n158 ? 1'b1 : 1'b0;
assign n2671 = /* LUT   18  9  4 */ n1287 ? 1'b1 : 1'b0;
assign n1364 = /* LUT   18 18  5 */ n718 ? n1118 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1118 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2673 = /* LUT    6 11  3 */ n115 ? n70 ? 1'b0 : n81 ? 1'b0 : 1'b1 : n70 ? n81 ? 1'b0 : 1'b1 : 1'b0;
assign n2674 = /* LUT   14 10  1 */ n414 ? 1'b1 : 1'b0;
assign n1478 = /* LUT   19 17  4 */ n1112 ? n709 ? n930 ? 1'b0 : 1'b1 : n993 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n993 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2676 = /* LUT   22 21  7 */ n218 ? 1'b1 : 1'b0;
assign n2677 = /* LUT    5 17  2 */ n87 ? n17 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n17 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2678 = /* LUT   24 13  0 */ n44 ? 1'b1 : 1'b0;
assign n2679 = /* LUT   21 14  1 */ n1431 ? n1648 ? n575 ? 1'b1 : 1'b0 : n1545 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1648 ? 1'b0 : n1545 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2680 = /* LUT    9 16  2 */ n235 ? n239 ? n236 ? n237 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2681 = /* LUT   14 20  6 */ n867 ? n190 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n190 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2682 = /* LUT   14  9  5 */ n751 ? n666 ? 1'b1 : n195 ? 1'b1 : 1'b0 : n666 ? n195 ? 1'b0 : 1'b1 : 1'b0;
assign n2683 = /* LUT   17 20  1 */ n397 ? 1'b0 : 1'b1;
assign n2684 = /* LUT   19 18  6 */ n1359 ? n687 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n687 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2685 = /* LUT   10 10  2 */ n288 ? 1'b1 : 1'b0;
assign n2686 = /* LUT   23 15  6 */ n140 ? 1'b1 : 1'b0;
assign n2687 = /* LUT   21 16  0 */ n44 ? 1'b1 : 1'b0;
assign n2688 = /* LUT   15 10  7 */ n919 ? 1'b1 : 1'b0;
assign n2689 = /* LUT   12  9  3 */ n295 ? 1'b0 : n286 ? 1'b0 : n296 ? 1'b0 : n294 ? 1'b0 : 1'b1;
assign n1399 = /* LUT   18 22  2 */ n731 ? n1127 ? 1'b1 : 1'b0 : 1'b0;
assign n2690 = /* LUT   11 19  2 */ n259 ? 1'b0 : 1'b1;
assign n2691 = /* LUT    9 12  4 */ n66 ? 1'b0 : n110 ? 1'b1 : 1'b0;
assign n2692 = /* LUT   13 17  0 */ n345 ? 1'b0 : n184 ? 1'b0 : n185 ? 1'b0 : n494 ? 1'b0 : 1'b1;
assign n2693 = /* LUT   18 21  4 */ n731 ? n885 ? n1127 ? n57 ? 1'b1 : 1'b0 : 1'b1 : n1127 ? n57 ? 1'b1 : 1'b0 : 1'b0 : n885 ? 1'b1 : 1'b0;
assign n2694 = /* LUT   19 14  5 */ n1318 ? n1452 ? n1059 ? n709 ? 1'b0 : 1'b1 : 1'b1 : n1059 ? 1'b0 : 1'b1 : n1452 ? n1059 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n1059 ? 1'b0 : n709 ? 1'b1 : 1'b0;
assign n2695 = /* LUT   22 20  4 */ n1678 ? n1741 ? n709 ? 1'b1 : 1'b0 : n709 ? n1234 ? 1'b1 : 1'b0 : 1'b1 : n1741 ? 1'b0 : n709 ? n1234 ? 1'b1 : 1'b0 : 1'b1;
assign n2696 = /* LUT   10 14  7 */ n208 ? 1'b0 : n211 ? 1'b0 : n209 ? 1'b0 : n210 ? 1'b0 : 1'b1;
assign n2697 = /* LUT    5 18  3 */ n96 ? n55 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n55 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2698 = /* LUT   16 24  5 */ io_4_33_0 ? 1'b1 : 1'b0;
assign n2699 = /* LUT    9 17  1 */ n159 ? 1'b1 : 1'b0;
assign n2700 = /* LUT   14 23  7 */ n212 ? 1'b1 : 1'b0;
assign n2701 = /* LUT   20 12  6 */ n140 ? 1'b1 : 1'b0;
assign n2702 = /* LUT   19 19  5 */ n140 ? 1'b1 : 1'b0;
assign n2703 = /* LUT   10 13  3 */ n308 ? n208 ? 1'b0 : n120 ? 1'b0 : 1'b1 : n208 ? n120 ? 1'b0 : 1'b1 : 1'b0;
assign n2704 = /* LUT   23 12  7 */ n218 ? 1'b1 : 1'b0;
assign n2705 = /* LUT   21 17  3 */ n35 ? 1'b1 : 1'b0;
assign n2706 = /* LUT   15 11  4 */ n278 ? 1'b1 : 1'b0;
assign n2707 = /* LUT   18 25  3 */ n1419 ? n575 ? n1420 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n1420 ? 1'b1 : 1'b0 : 1'b0;
assign n2708 = /* LUT   20 15  0 */ n180 ? 1'b0 : n932 ? 1'b0 : n244 ? n238 ? 1'b1 : 1'b0 : 1'b0;
assign n2709 = /* LUT   11 16  3 */ n355 ? 1'b1 : 1'b0;
assign n2710 = /* LUT   16  9  0 */ n159 ? 1'b1 : 1'b0;
assign n2711 = /* LUT   13 18  1 */ n256 ? 1'b0 : 1'b1;
assign n2712 = /* LUT   15 20  2 */ n720 ? 1'b0 : 1'b1;
assign n2713 = /* LUT   18 20  7 */ n1128 ? n709 ? n930 ? 1'b0 : 1'b1 : n1275 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1275 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2714 = /* LUT   16  7  3 */ n1050 ? n903 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n903 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n1465 = /* LUT   19 15  6 */ n1208 ? n1460 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1460 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n2716 = /* LUT   22 23  5 */ n158 ? 1'b1 : 1'b0;
assign n2717 = /* LUT   15 26  1 */ n1045 ? n899 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n899 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2718 = /* LUT    9 18  0 */ n35 ? 1'b1 : 1'b0;
assign n2719 = /* LUT   12 12  1 */ n427 ? 1'b1 : 1'b0;
assign n2720 = /* LUT   14 22  0 */ n159 ? 1'b1 : 1'b0;
assign n2721 = /* LUT   17 22  3 */ n981 ? 1'b0 : 1'b1;
assign n2722 = /* LUT   14 11  7 */ n663 ? 1'b1 : 1'b0;
assign n2723 = /* LUT   19 16  4 */ n35 ? 1'b1 : 1'b0;
assign n2727 = /* LUT   21 18  2 */ n44 ? 1'b1 : 1'b0;
assign n2728 = /* LUT   12 15  5 */ n488 ? 1'b0 : 1'b1;
assign n2729 = /* LUT   15  7  4 */ n905 ? 1'b0 : n907 ? n902 ? 1'b1 : 1'b0 : 1'b0;
assign n1569 = /* LUT   20 14  3 */ n1237 ? n709 ? n930 ? 1'b0 : 1'b1 : n1457 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1457 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2731 = /* LUT   23 20  0 */ n159 ? 1'b1 : 1'b0;
assign n2732 = /* LUT   13 19  6 */ n188 ? 1'b0 : 1'b1;
assign n2733 = /* LUT   18 23  6 */ n731 ? n896 ? n1127 ? n58 ? 1'b1 : 1'b0 : 1'b1 : n1127 ? n58 ? 1'b1 : 1'b0 : 1'b0 : n896 ? 1'b1 : 1'b0;
assign n2734 = /* LUT   14 18  5 */ n832 ? n345 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n345 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2735 = /* LUT   14  7  2 */ n742 ? n648 ? 1'b0 : n734 ? 1'b0 : 1'b1 : n648 ? n734 ? 1'b0 : 1'b1 : 1'b0;
assign n2736 = /* LUT   19 12  7 */ n180 ? n1435 ? 1'b1 : 1'b0 : 1'b0;
assign n2737 = /* LUT   12 19  0 */ n159 ? 1'b1 : 1'b0;
assign n2738 = /* LUT   14 17  1 */ n397 ? 1'b0 : n190 ? 1'b0 : n189 ? 1'b0 : n396 ? 1'b0 : 1'b1;
assign n2739 = /* LUT   17 12  5 */ n439 ? n1159 ? 1'b1 : n575 ? 1'b1 : 1'b0 : n1159 ? n575 ? 1'b0 : 1'b1 : 1'b0;
assign n2740 = /* LUT   17 23  4 */ n877 ? 1'b0 : 1'b1;
assign n2741 = /* LUT   10 15  1 */ n332 ? n220 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n220 ? 1'b1 : 1'b0;
assign n1684 = /* LUT   21 19  5 */ n1601 ? n1683 ? n705 ? 1'b0 : 1'b1 : 1'b0 : n1552 ? 1'b1 : n705 ? 1'b1 : 1'b0;
assign n2745 = /* LUT   18 14  6 */ n712 ? n1190 ? 1'b1 : 1'b0 : n960 ? 1'b1 : 1'b0;
assign n2746 = /* LUT   15  9  2 */ n915 ? 1'b1 : 1'b0;
assign n2747 = /* LUT   12 14  6 */ n490 ? 1'b0 : 1'b1;
assign n2748 = /* LUT   20 13  2 */ n1436 ? n1557 ? n930 ? 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? 1'b0 : 1'b1 : n1557 ? n930 ? n709 ? 1'b1 : 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? n709 ? 1'b1 : 1'b0 : 1'b1;
assign n2749 = /* LUT   10 17  5 */ n364 ? n228 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n228 ? 1'b1 : 1'b0;
assign n2750 = /* LUT    9 15  1 */ n219 ? n228 ? n213 ? n227 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2751 = /* LUT   13 20  7 */ n526 ? 1'b0 : 1'b1;
assign n1312 = /* LUT   18 13  0 */ n1184 ? n705 ? n1183 ? 1'b0 : 1'b1 : n1183 ? 1'b1 : n1311 ? 1'b1 : 1'b0 : n705 ? n1183 ? 1'b0 : 1'b1 : n1183 ? 1'b0 : n1311 ? 1'b1 : 1'b0;
assign n2753 = /* LUT   20 19  1 */ n212 ? 1'b1 : 1'b0;
assign n2754 = /* LUT   14 13  4 */ n35 ? 1'b1 : 1'b0;
assign n2757 = /* LUT   19 13  0 */ n159 ? 1'b1 : 1'b0;
assign n2758 = /* LUT   22 17  3 */ n1617 ? n1731 ? n1584 ? n709 ? 1'b1 : 1'b0 : 1'b0 : 1'b1 : n1731 ? n1584 ? n709 ? 1'b1 : 1'b0 : 1'b0 : n709 ? 1'b0 : 1'b1;
assign n2759 = /* LUT   15 24  3 */ n1029 ? n887 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n887 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2760 = /* LUT   21 23  2 */ n35 ? 1'b1 : 1'b0;
assign n2761 = /* LUT   15 13  7 */ n140 ? n770 ? 1'b0 : 1'b1 : 1'b0;
assign n2762 = /* LUT   12 18  3 */ n612 ? n487 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n487 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2763 = /* LUT   14 16  2 */ n700 ? 1'b1 : 1'b0;
assign n1189 = /* LUT   17 13  6 */ n952 ? n1180 ? 1'b1 : n1176 ? 1'b1 : 1'b0 : n1180 ? 1'b0 : n1176 ? 1'b1 : 1'b0;
assign n1214 = /* LUT   17 16  5 */ n1100 ? n1213 ? n709 ? n930 ? 1'b0 : 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n930 ? 1'b1 : 1'b0 : n1213 ? n930 ? 1'b0 : 1'b1 : n709 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2766 = /* LUT   21 20  4 */ n35 ? 1'b1 : 1'b0;
assign n2769 = /* LUT   15 14  3 */ n591 ? n770 ? n776 ? 1'b0 : n771 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2770 = /* LUT   18 17  7 */ n1351 ? n1113 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1113 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2771 = /* LUT   12 13  7 */ n218 ? 1'b1 : 1'b0;
assign n2772 = /* LUT   10 16  6 */ n351 ? n236 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n236 ? 1'b1 : 1'b0;
assign n2773 = /* LUT   18 12  3 */ n42 ? 1'b1 : 1'b0;
assign n2774 = /* LUT   20 18  2 */ n782 ? n159 ? n703 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2775 = /* LUT   19 10  1 */ n212 ? 1'b1 : 1'b0;
assign n2776 = /* LUT   22 16  0 */ n42 ? 1'b1 : 1'b0;
assign n2777 = /* LUT   15 25  4 */ n1039 ? n541 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n541 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2778 = /* LUT   12 17  2 */ n598 ? n470 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n470 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2779 = /* LUT   14 19  3 */ n847 ? n514 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n514 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2780 = /* LUT   17 14  7 */ n968 ? n1198 ? n575 ? 1'b1 : 1'b0 : n791 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1198 ? 1'b0 : n791 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2781 = /* LUT   19 24  0 */ n1525 ? n1405 ? 1'b0 : n1501 ? 1'b0 : 1'b1 : n1405 ? n1501 ? 1'b0 : 1'b1 : 1'b0;
assign n2782 = /* LUT   17 17  6 */ n1110 ? n1221 ? n1180 ? 1'b0 : 1'b1 : 1'b0 : n1221 ? n705 ? n1180 ? 1'b0 : 1'b1 : 1'b1 : 1'b0;
assign n2783 = /* LUT   21 21  7 */ n1149 ? n709 ? n930 ? 1'b0 : 1'b1 : n1616 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1616 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2784 = /* LUT   15 15  0 */ n159 ? 1'b1 : 1'b0;
assign n2785 = /* LUT   18 16  4 */ n1345 ? n712 ? n1180 ? 1'b0 : 1'b1 : 1'b0 : n712 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n2786 = /* LUT   10 19  7 */ n218 ? 1'b1 : 1'b0;
assign n2787 = /* LUT   13 11  2 */ n566 ? n559 ? 1'b0 : io_33_1_1 ? 1'b1 : n561 ? 1'b0 : 1'b1 : n559 ? io_33_1_1 ? 1'b1 : n561 ? 1'b0 : 1'b1 : 1'b0;
assign n2788 = /* LUT   13 22  5 */ n403 ? 1'b0 : 1'b1;
assign n1333 = /* LUT   18 15  2 */ n1104 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1200 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1200 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2790 = /* LUT    6 12  2 */ n70 ? n69 ? 1'b1 : n67 ? 1'b1 : n68 ? 1'b0 : 1'b1 : 1'b1;
assign n2791 = /* LUT   20 17  3 */ n212 ? 1'b1 : 1'b0;
assign n2792 = /* LUT   14 15  6 */ n798 ? n771 ? 1'b1 : 1'b0 : 1'b0;
assign n2793 = /* LUT   19 11  2 */ n44 ? 1'b1 : 1'b0;
assign n2794 = /* LUT   22 19  1 */ n35 ? 1'b1 : 1'b0;
assign n2795 = /* LUT   12 16  5 */ n481 ? io_0_27_1 ? n341 ? 1'b1 : n340 ? 1'b1 : 1'b0 : n341 ? 1'b1 : 1'b0 : n341 ? 1'b1 : 1'b0;
assign n1205 = /* LUT   17 15  0 */ n1088 ? n575 ? n1180 ? 1'b0 : 1'b1 : n804 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n804 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2799 = /* LUT   22 13  5 */ n35 ? 1'b1 : 1'b0;
assign n2800 = /* LUT   15 12  1 */ n358 ? n691 ? 1'b1 : n591 ? n934 ? 1'b1 : 1'b0 : 1'b1 : n691 ? n591 ? 1'b1 : 1'b0 : n591 ? n934 ? 1'b1 : 1'b0 : 1'b0;
assign n2801 = /* LUT   18 19  5 */ n1374 ? n1228 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1228 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2802 = /* LUT   11 22  1 */ n212 ? 1'b1 : 1'b0;
assign n2803 = /* LUT   16 15  2 */ n59 ? n802 ? n244 ? 1'b0 : n948 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2804 = /* LUT   10 18  0 */ n365 ? n239 ? 1'b0 : 1'b1 : n239 ? 1'b1 : 1'b0;
assign n2805 = /* LUT   13 12  3 */ n680 ? n567 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n567 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2806 = /* LUT   15 18  0 */ n159 ? 1'b1 : 1'b0;
assign n2807 = /* LUT   20 16  4 */ n35 ? 1'b1 : 1'b0;
assign n2808 = /* LUT   12 20  2 */ n44 ? 1'b1 : 1'b0;
assign n2810 = /* LUT   17 11  5 */ n1166 ? n927 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n927 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2811 = /* LUT   19  8  3 */ n1423 ? 1'b1 : 1'b0;
assign n2812 = /* LUT   23 14  0 */ n159 ? 1'b1 : 1'b0;
assign n2813 = /* LUT   24 17  0 */ n159 ? 1'b1 : 1'b0;
assign n2814 = /* LUT   21 10  1 */ n1424 ? n1628 ? n1623 ? n1540 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2815 = /* LUT   12 10  7 */ n152 ? n554 ? 1'b1 : 1'b0 : n548 ? 1'b1 : 1'b0;
assign n2818 = /* LUT   17  8  1 */ n1157 ? 1'b1 : 1'b0;
assign n2819 = /* LUT   16 16  0 */ n159 ? 1'b1 : 1'b0;
assign n2820 = /* LUT   22 12  6 */ n140 ? 1'b1 : 1'b0;
assign n2821 = /* LUT   13 16  6 */ n159 ? 1'b1 : 1'b0;
assign n137  = /* LUT    7 12  6 */ n66 ? 1'b0 : n107 ? 1'b1 : n110 ? 1'b1 : 1'b0;
assign n2822 = /* LUT   18 18  2 */ n1239 ? n1363 ? n709 ? 1'b1 : 1'b0 : 1'b0 : n1222 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n2823 = /* LUT   20 20  1 */ n212 ? 1'b1 : 1'b0;
assign n2824 = /* LUT   23 18  2 */ n42 ? 1'b1 : 1'b0;
assign n2825 = /* LUT   16 14  1 */ n780 ? n778 ? n935 ? n943 ? 1'b0 : 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2826 = /* LUT    5 17  7 */ n92 ? n27 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n27 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2827 = /* LUT   13 13  0 */ n569 ? 1'b0 : n559 ? n557 ? 1'b1 : 1'b0 : 1'b0;
assign n2828 = /* LUT   15 19  3 */ n42 ? 1'b1 : 1'b0;
assign n2829 = /* LUT   20 23  5 */ n44 ? 1'b1 : 1'b0;
assign n2830 = /* LUT   14  9  0 */ n667 ? n748 ? 1'b1 : n152 ? 1'b1 : 1'b0 : n748 ? n152 ? 1'b0 : 1'b1 : 1'b0;
assign n2831 = /* LUT   17 20  4 */ n189 ? 1'b0 : 1'b1;
assign n2832 = /* LUT   23 15  3 */ n42 ? 1'b1 : 1'b0;
assign n2833 = /* LUT   21 16  7 */ n1581 ? n1666 ? n709 ? n1572 ? 1'b0 : 1'b1 : 1'b1 : n709 ? n1572 ? 1'b0 : 1'b1 : n1572 ? 1'b1 : 1'b0 : n1666 ? n1572 ? 1'b0 : 1'b1 : n709 ? n1572 ? 1'b0 : 1'b1 : 1'b0;
assign n2834 = /* LUT   21 11  6 */ n140 ? 1'b1 : 1'b0;
assign n2835 = /* LUT   18 22  7 */ n272 ? io_0_25_1 ? n1021 ? n1025 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0;
assign n2838 = /* LUT   10  9  3 */ n136 ? 1'b1 : 1'b0;
assign n2839 = /* LUT   22 15  7 */ n59 ? n525 ? 1'b0 : n244 ? n238 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2840 = /* LUT   13 17  5 */ n385 ? 1'b0 : n184 ? 1'b0 : n183 ? 1'b0 : n185 ? 1'b0 : 1'b1;
assign n2841 = /* LUT   18 21  3 */ n17 ? n1127 ? n731 ? 1'b1 : n884 ? 1'b1 : 1'b0 : n884 ? 1'b1 : 1'b0 : n1127 ? n731 ? 1'b0 : n884 ? 1'b1 : 1'b0 : n884 ? 1'b1 : 1'b0;
assign n2842 = /* LUT   20 11  0 */ n212 ? 1'b1 : 1'b0;
assign n2843 = /* LUT   23 19  1 */ n1710 ? n575 ? n1744 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n1744 ? 1'b1 : 1'b0 : 1'b0;
assign n2844 = /* LUT   11 20  3 */ n250 ? 1'b0 : 1'b1;
assign n2845 = /* LUT   16 13  0 */ n590 ? n244 ? n932 ? 1'b0 : n180 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2846 = /* LUT    5 18  6 */ n99 ? n58 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n58 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2847 = /* LUT   10 20  2 */ n35 ? 1'b1 : 1'b0;
assign n2848 = /* LUT   15 16  2 */ n590 ? n59 ? 1'b0 : n244 ? n525 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n1658 = /* LUT   21 15  3 */ n1576 ? n1544 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1544 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2850 = /* LUT   20 25  7 */ n218 ? 1'b1 : 1'b0;
assign n2851 = /* LUT   20 22  6 */ n731 ? n1501 ? n1127 ? io_11_33_1 ? 1'b0 : 1'b1 : 1'b0 : n1127 ? io_11_33_1 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2854 = /* LUT   23 12  2 */ n44 ? 1'b1 : 1'b0;
assign n2855 = /* LUT    7 10  7 */ n75 ? n136 ? 1'b1 : 1'b0 : 1'b0;
assign n2856 = /* LUT   21 17  4 */ n1588 ? n575 ? n1598 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n1598 ? 1'b1 : 1'b0 : 1'b0;
assign n2857 = /* LUT   21 12  7 */ n218 ? 1'b1 : 1'b0;
assign n2858 = /* LUT   18 25  6 */ n1416 ? n575 ? n1415 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n1415 ? 1'b1 : 1'b0 : 1'b0;
assign n2859 = /* LUT   12 21  6 */ n522 ? 1'b0 : 1'b1;
assign n2860 = /* LUT   22 14  0 */ n159 ? 1'b1 : 1'b0;
assign n2861 = /* LUT   13 18  4 */ n183 ? 1'b0 : 1'b1;
assign n1385 = /* LUT   18 20  0 */ n1248 ? n1384 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1384 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2863 = /* LUT   20 10  3 */ n1425 ? 1'b0 : 1'b1;
assign n2864 = /* LUT   23 16  0 */ n159 ? 1'b1 : 1'b0;
assign n2865 = /* LUT   11 14  5 */ n455 ? n436 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n436 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n2866 = /* LUT   16 12  7 */ n776 ? 1'b1 : n1072 ? 1'b1 : n180 ? 1'b1 : n244 ? 1'b0 : 1'b1;
assign n2867 = /* LUT    5 19  1 */ n102 ? n61 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n61 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2868 = /* LUT   22 24  1 */ n218 ? 1'b1 : 1'b0;
assign n2869 = /* LUT   15 17  5 */ n158 ? 1'b1 : 1'b0;
assign n2870 = /* LUT   12 12  6 */ n423 ? 1'b1 : 1'b0;
assign n2871 = /* LUT   20 21  7 */ n140 ? 1'b1 : 1'b0;
assign n2872 = /* LUT   17 22  6 */ n861 ? 1'b0 : 1'b1;
assign n2873 = /* LUT   14 11  2 */ n658 ? 1'b1 : 1'b0;
assign n2874 = /* LUT   22 10  5 */ n1705 ? 1'b1 : 1'b0;
assign n2875 = /* LUT   21 18  5 */ n42 ? 1'b1 : 1'b0;
assign n2876 = /* LUT   21 13  4 */ n212 ? 1'b1 : 1'b0;
assign n2877 = /* LUT   12 15  0 */ n484 ? 1'b0 : 1'b1;
assign n906  = /* LUT   15  7  1 */ n738 ? n647 ? n648 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2878 = /* LUT   18 24  5 */ n1271 ? n1414 ? n709 ? 1'b1 : 1'b0 : n1277 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1414 ? 1'b0 : n1277 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n2879 = /* LUT   11 17  1 */ n342 ? 1'b0 : io_0_25_1 ? 1'b1 : 1'b0;
assign n2880 = /* LUT   13 19  3 */ n514 ? 1'b0 : 1'b1;
assign n2881 = /* LUT   15 21  2 */ n998 ? 1'b0 : 1'b1;
assign n2882 = /* LUT   18 23  1 */ n50 ? n1127 ? n731 ? 1'b1 : n890 ? 1'b1 : 1'b0 : n890 ? 1'b1 : 1'b0 : n1127 ? n731 ? 1'b0 : n890 ? 1'b1 : 1'b0 : n890 ? 1'b1 : 1'b0;
assign n2883 = /* LUT   23 17  7 */ n1743 ? n1747 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1747 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2884 = /* LUT   11 15  6 */ n479 ? n301 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n301 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n2885 = /* LUT   14  7  5 */ n745 ? n651 ? 1'b0 : 1'b1 : n651 ? 1'b1 : 1'b0;
assign n2886 = /* LUT   11 18  5 */ n508 ? 1'b0 : 1'b1;
assign n2887 = /* LUT   16 11  6 */ n140 ? 1'b1 : 1'b0;
assign n2890 = /* LUT   18  9  0 */ n135 ? 1'b1 : 1'b0;
assign n2891 = /* LUT   12 19  7 */ n218 ? 1'b1 : 1'b0;
assign n2892 = /* LUT    6 11  7 */ n119 ? n81 ? 1'b0 : n74 ? 1'b0 : 1'b1 : n81 ? 1'b0 : n74 ? 1'b1 : 1'b0;
assign n2893 = /* LUT   17 23  1 */ n992 ? 1'b0 : 1'b1;
assign n1476 = /* LUT   19 17  0 */ n1346 ? n709 ? n1456 ? 1'b1 : 1'b0 : 1'b0 : n709 ? n959 ? 1'b1 : 1'b0 : 1'b1;
assign n2895 = /* LUT   22 21  3 */ n42 ? 1'b1 : 1'b0;
assign n2896 = /* LUT    7  8  5 */ n65 ? 1'b1 : 1'b0;
assign n2897 = /* LUT   21 19  2 */ n1679 ? n1681 ? n595 ? 1'b0 : n705 ? 1'b0 : 1'b1 : n595 ? 1'b0 : 1'b1 : n1681 ? n595 ? n705 ? 1'b1 : 1'b0 : n705 ? 1'b0 : 1'b1 : n595 ? n705 ? 1'b1 : 1'b0 : 1'b1;
assign n2898 = /* LUT   21 14  5 */ n212 ? 1'b1 : 1'b0;
assign n2899 = /* LUT   12 14  3 */ n471 ? 1'b0 : 1'b1;
assign n2900 = /* LUT   14 20  2 */ n863 ? n528 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n528 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2903 = /* LUT   16 23  5 */ n468 ? 1'b1 : 1'b0;
assign n2904 = /* LUT   13 20  2 */ n528 ? 1'b0 : 1'b1;
assign n2905 = /* LUT   20 19  4 */ n35 ? 1'b1 : 1'b0;
assign n2906 = /* LUT   11 12  7 */ n428 ? 1'b1 : 1'b0;
assign n2909 = /* LUT   11 19  6 */ n263 ? 1'b0 : 1'b1;
assign n2910 = /* LUT   16 10  5 */ n1047 ? 1'b1 : 1'b0;
assign n2911 = /* LUT   15 24  6 */ n1032 ? n890 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n890 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2912 = /* LUT   12 18  4 */ n613 ? n499 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n499 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2913 = /* LUT   17 16  0 */ n1101 ? n575 ? 1'b1 : n1210 ? 1'b1 : 1'b0 : n575 ? 1'b0 : n1210 ? 1'b1 : 1'b0;
assign n1450 = /* LUT   19 14  1 */ n1449 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1292 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1292 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2915 = /* LUT   22 20  0 */ n1614 ? n709 ? n1685 ? 1'b1 : 1'b0 : 1'b0 : n709 ? n1688 ? 1'b1 : 1'b0 : 1'b1;
assign n2916 = /* LUT   10 14  3 */ io_0_25_1 ? n322 ? 1'b1 : 1'b0 : 1'b0;
assign n2917 = /* LUT   16 24  1 */ io_6_33_1 ? 1'b1 : 1'b0;
assign n2918 = /* LUT   21 20  3 */ n42 ? 1'b1 : 1'b0;
assign n2919 = /* LUT    9 17  5 */ n212 ? 1'b1 : 1'b0;
assign n2920 = /* LUT   12 13  2 */ n44 ? 1'b1 : 1'b0;
assign n2921 = /* LUT   20 12  2 */ n44 ? 1'b1 : 1'b0;
assign n2922 = /* LUT   10 13  7 */ n312 ? n120 ? 1'b0 : n211 ? 1'b0 : 1'b1 : n120 ? 1'b0 : n211 ? 1'b1 : 1'b0;
assign n2923 = /* LUT   15 11  0 */ n931 ? 1'b1 : 1'b0;
assign n1578 = /* LUT   20 15  4 */ n1302 ? n180 ? 1'b0 : 1'b1 : 1'b0;
assign n2924 = /* LUT   11 13  0 */ n44 ? 1'b1 : 1'b0;
assign n2925 = /* LUT   11 16  7 */ n51 ? n343 ? 1'b0 : n358 ? 1'b1 : 1'b0 : n343 ? n169 ? 1'b0 : 1'b1 : n169 ? n358 ? 1'b1 : 1'b0 : 1'b1;
assign n656  = /* LUT   13  7  2 */ n647 ? n645 ? 1'b1 : 1'b0 : n655 ? 1'b1 : 1'b0;
assign n2927 = /* LUT   15 25  1 */ n1036 ? n892 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n892 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n2928 = /* LUT   18 11  2 */ n44 ? 1'b1 : 1'b0;
assign n2929 = /* LUT   15 20  6 */ n841 ? 1'b0 : 1'b1;
assign n2930 = /* LUT   12 17  5 */ n601 ? n473 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n473 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n2931 = /* LUT   17 17  3 */ n986 ? n923 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n923 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2932 = /* LUT   19 15  2 */ n1327 ? n1463 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1463 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2933 = /* LUT   22 23  1 */ n212 ? 1'b1 : 1'b0;
assign n1695 = /* LUT   21 21  0 */ n1613 ? n1493 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1493 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2935 = /* LUT   14 22  4 */ n140 ? 1'b1 : 1'b0;
assign n2936 = /* LUT   11  9  5 */ n279 ? n278 ? 1'b1 : n150 ? 1'b1 : 1'b0 : n278 ? n150 ? n65 ? 1'b1 : 1'b0 : 1'b1 : 1'b0;
assign n2937 = /* LUT   16 21  7 */ n212 ? 1'b1 : 1'b0;
assign n2938 = /* LUT   13 22  0 */ n145 ? 1'b0 : 1'b1;
assign n2940 = /* LUT   15  8  1 */ n545 ? n912 ? 1'b1 : n647 ? 1'b1 : 1'b0 : n912 ? n647 ? 1'b0 : 1'b1 : 1'b0;
assign n2941 = /* LUT   20 17  6 */ n1474 ? n1226 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1226 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2942 = /* LUT   23 20  4 */ n35 ? 1'b1 : 1'b0;
assign n2943 = /* LUT   11 10  1 */ n293 ? n412 ? n154 ? n284 ? 1'b1 : 1'b0 : 1'b1 : 1'b1 : n412 ? n154 ? n284 ? 1'b1 : 1'b0 : 1'b1 : 1'b0;
assign n2944 = /* LUT    9 14  2 */ n160 ? n84 ? n165 ? n161 ? 1'b0 : 1'b1 : 1'b1 : n165 ? n161 ? 1'b1 : 1'b0 : 1'b0 : n84 ? 1'b1 : 1'b0;
assign n2945 = /* LUT   14 18  1 */ n828 ? n256 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n256 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n2948 = /* LUT   19 12  3 */ n590 ? n802 ? n244 ? n59 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2949 = /* LUT   21 22  1 */ n1615 ? n1605 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1605 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2950 = /* LUT   14 17  5 */ n712 ? n818 ? 1'b1 : 1'b0 : n795 ? 1'b1 : 1'b0;
assign n1182 = /* LUT   17 12  1 */ n942 ? n941 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n941 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n2952 = /* LUT   11 22  4 */ n35 ? 1'b1 : 1'b0;
assign n2953 = /* LUT   10 15  5 */ n336 ? n224 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n224 ? 1'b1 : 1'b0;
assign n2954 = /* LUT   16 20  0 */ n1025 ? io_11_33_1 ? io_0_25_1 ? 1'b1 : n994 ? 1'b1 : 1'b0 : io_0_25_1 ? 1'b0 : n994 ? 1'b1 : 1'b0 : n994 ? 1'b1 : 1'b0;
assign n2955 = /* LUT   21 24  0 */ n35 ? 1'b1 : 1'b0;
assign n2956 = /* LUT   15 18  7 */ n218 ? 1'b1 : 1'b0;
assign n1325 = /* LUT   18 14  2 */ n1323 ? n709 ? n930 ? 1'b0 : 1'b1 : n1306 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1306 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2958 = /* LUT   20 16  1 */ n212 ? 1'b1 : 1'b0;
assign n2959 = /* LUT   12 20  7 */ n218 ? 1'b1 : 1'b0;
assign n2960 = /* LUT   20 13  6 */ n1296 ? n925 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n925 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2961 = /* LUT   11 11  2 */ n417 ? n294 ? 1'b0 : n282 ? 1'b0 : 1'b1 : n294 ? n282 ? 1'b0 : 1'b1 : 1'b0;
assign n2962 = /* LUT   22 18  3 */ n1728 ? n709 ? n930 ? 1'b0 : 1'b1 : n1356 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1356 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n2963 = /* LUT   10 17  1 */ n360 ? n240 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n240 ? 1'b1 : 1'b0;
assign n230  = /* LUT    9 15  5 */ n159 ? 1'b0 : n140 ? 1'b0 : 1'b1;
assign n2965 = /* LUT   13  9  0 */ n14 ? 1'b1 : 1'b0;
assign n1629 = /* LUT   21 10  4 */ n1535 ? n1294 ? n1624 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2967 = /* LUT   18 13  4 */ n1195 ? n1314 ? n595 ? 1'b0 : n705 ? 1'b0 : 1'b1 : n595 ? 1'b0 : 1'b1 : n1314 ? n595 ? n705 ? 1'b1 : 1'b0 : n705 ? 1'b0 : 1'b1 : n595 ? n705 ? 1'b1 : 1'b0 : 1'b1;
assign n2970 = /* LUT   14 13  0 */ n159 ? 1'b1 : 1'b0;
assign n2971 = /* LUT   19 22  5 */ n1515 ? n1394 ? 1'b0 : n1258 ? 1'b0 : 1'b1 : n1394 ? n1258 ? 1'b0 : 1'b1 : 1'b0;
assign n2972 = /* LUT   19 13  4 */ n1307 ? n217 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n217 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n2973 = /* LUT   16 16  5 */ n158 ? 1'b1 : 1'b0;
assign n2974 = /* LUT    7 12  1 */ n14 ? 1'b0 : n125 ? 1'b1 : 1'b0;
assign n2975 = /* LUT   15 13  3 */ n591 ? n775 ? n782 ? n777 ? 1'b0 : 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n2976 = /* LUT   20 20  6 */ n140 ? 1'b1 : 1'b0;
assign n2977 = /* LUT   14 16  6 */ n696 ? io_33_1_1 ? 1'b1 : n320 ? 1'b1 : io_0_25_1 ? 1'b0 : 1'b1 : io_33_1_1 ? n320 ? 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n320 ? 1'b1 : 1'b0;
assign n2978 = /* LUT   17 13  2 */ n1073 ? n1187 ? n575 ? 1'b1 : 1'b0 : n1085 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1187 ? 1'b0 : n1085 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n2979 = /* LUT   16 19  1 */ n42 ? 1'b1 : 1'b0;
assign n2980 = /* LUT   15 19  4 */ n35 ? 1'b1 : 1'b0;
assign n2981 = /* LUT   18 17  3 */ n218 ? 1'b1 : 1'b0;
assign n2982 = /* LUT   15 14  7 */ n591 ? n957 ? n779 ? 1'b0 : n689 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2983 = /* LUT   20 23  0 */ n1523 ? n692 ? n1522 ? n1524 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n2984 = /* LUT   10 16  2 */ n347 ? n232 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n232 ? 1'b1 : 1'b0;
assign n2985 = /* LUT   13 10  1 */ n661 ? 1'b1 : 1'b0;
assign n2986 = /* LUT   21 11  3 */ n42 ? 1'b1 : 1'b0;
assign n2987 = /* LUT   18 12  7 */ n218 ? 1'b1 : 1'b0;
assign n2990 = /* LUT   14 12  3 */ n767 ? n768 ? 1'b1 : n151 ? 1'b1 : 1'b0 : n768 ? n151 ? 1'b0 : 1'b1 : 1'b0;
assign n2991 = /* LUT   19 23  6 */ n1025 ? io_0_25_1 ? n272 ? n1404 ? 1'b1 : 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n2992 = /* LUT   19 10  5 */ n158 ? 1'b1 : 1'b0;
assign n2993 = /* LUT   22 16  4 */ n686 ? n1723 ? 1'b1 : n575 ? 1'b1 : 1'b0 : n1723 ? n575 ? 1'b0 : 1'b1 : 1'b0;
assign n2994 = /* LUT   14 19  7 */ n851 ? n513 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n513 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n1197 = /* LUT   17 14  3 */ n1082 ? n575 ? n1180 ? 1'b0 : 1'b1 : n970 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n970 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n2996 = /* LUT   19 24  4 */ n1529 ? n1409 ? 1'b0 : n1501 ? 1'b0 : 1'b1 : n1409 ? n1501 ? 1'b0 : 1'b1 : 1'b0;
assign n2997 = /* LUT   11 20  6 */ n253 ? 1'b0 : 1'b1;
assign n2998 = /* LUT   16 18  2 */ n44 ? 1'b1 : 1'b0;
assign n2999 = /* LUT   15 16  5 */ n141 ? n244 ? 1'b0 : n180 ? n59 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n3000 = /* LUT   15 15  4 */ n35 ? 1'b1 : 1'b0;
assign n1619 = /* LUT   20 22  3 */ n1392 ? n1395 ? 1'b1 : n1504 ? 1'b0 : 1'b1 : 1'b1;
assign n3007 = /* LUT   10 19  3 */ n42 ? 1'b1 : 1'b0;
assign n3008 = /* LUT   13 11  6 */ io_33_1_1 ? 1'b0 : 1'b1;
assign n3009 = /* LUT   21 12  2 */ n44 ? 1'b1 : 1'b0;
assign n3010 = /* LUT   18 15  6 */ n1201 ? n1335 ? n1106 ? n709 ? 1'b0 : 1'b1 : 1'b1 : n1106 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n1335 ? n1106 ? 1'b0 : 1'b1 : n1106 ? 1'b0 : n709 ? 1'b1 : 1'b0;
assign n3011 = /* LUT   12 21  1 */ n539 ? 1'b0 : 1'b1;
assign n3012 = /* LUT   19 20  7 */ n937 ? 1'b0 : n244 ? 1'b0 : n590 ? 1'b1 : 1'b0;
assign n3013 = /* LUT   19 11  6 */ n140 ? 1'b1 : 1'b0;
assign n3014 = /* LUT   22 19  5 */ n140 ? 1'b1 : 1'b0;
assign n3015 = /* LUT   17 15  4 */ n813 ? n1206 ? n575 ? n1153 ? 1'b1 : 1'b0 : 1'b0 : 1'b1 : n1206 ? n575 ? n1153 ? 1'b1 : 1'b0 : 1'b0 : n575 ? 1'b0 : 1'b1;
assign n3016 = /* LUT   16 17  3 */ n42 ? 1'b1 : 1'b0;
assign n3017 = /* LUT   22 13  1 */ n1548 ? n1713 ? n575 ? n1433 ? 1'b1 : 1'b0 : 1'b0 : 1'b1 : n1713 ? n575 ? n1433 ? 1'b1 : 1'b0 : 1'b0 : n575 ? 1'b0 : 1'b1;
assign n3018 = /* LUT   15 17  2 */ n44 ? 1'b1 : 1'b0;
assign n3019 = /* LUT   15 12  5 */ n740 ? io_33_1_1 ? 1'b1 : n571 ? 1'b1 : 1'b0 : io_33_1_1 ? 1'b0 : n571 ? 1'b1 : 1'b0;
assign n3020 = /* LUT   18 19  1 */ n140 ? 1'b1 : 1'b0;
assign n3021 = /* LUT   20 21  2 */ n1497 ? n1507 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1507 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3022 = /* LUT   17 25  0 */ n1274 ? 1'b0 : n374 ? n354 ? 1'b0 : n1109 ? 1'b1 : 1'b0 : n1109 ? 1'b1 : 1'b0;
assign n3023 = /* LUT   24 14  6 */ n140 ? 1'b1 : 1'b0;
assign n1643 = /* LUT   21 13  1 */ n1165 ? n1331 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1331 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n1168 = /* LUT   17 11  1 */ n1061 ? n570 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n570 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3026 = /* LUT   19 21  0 */ n1025 ? 1'b1 : n383 ? n641 ? n1011 ? 1'b1 : 1'b0 : 1'b1 : n641 ? n1011 ? 1'b1 : 1'b0 : 1'b0;
assign n498  = /* LUT   11 17  6 */ n183 ? n385 ? 1'b0 : 1'b1 : 1'b0;
assign n3028 = /* LUT   23 14  4 */ n35 ? 1'b1 : 1'b0;
assign n3029 = /* LUT   24 17  4 */ n35 ? 1'b1 : 1'b0;
assign n3030 = /* LUT   15 21  7 */ n1003 ? 1'b0 : 1'b1;
assign n3031 = /* LUT   12 10  3 */ n556 ? n553 ? 1'b1 : n195 ? 1'b0 : 1'b1 : n553 ? n195 ? 1'b1 : 1'b0 : 1'b0;
assign n3032 = /* LUT   17  8  5 */ n1155 ? 1'b1 : 1'b0;
assign n3033 = /* LUT   11 18  0 */ n503 ? 1'b0 : 1'b1;
assign n3035 = /* LUT   22 12  2 */ n44 ? 1'b1 : 1'b0;
assign n3036 = /* LUT   13 16  2 */ n35 ? 1'b1 : 1'b0;
assign n3039 = /* LUT   18  9  7 */ n1286 ? 1'b1 : 1'b0;
assign n1365 = /* LUT   18 18  6 */ n1225 ? n1364 ? n930 ? 1'b0 : n709 ? 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n1364 ? n930 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n930 ? n709 ? 1'b0 : 1'b1 : 1'b1;
assign n3041 = /* LUT    6 11  2 */ n114 ? n69 ? 1'b0 : n81 ? 1'b0 : 1'b1 : n69 ? n81 ? 1'b0 : 1'b1 : 1'b0;
assign n3042 = /* LUT   14 10  2 */ n673 ? 1'b1 : 1'b0;
assign n1479 = /* LUT   19 17  5 */ n1348 ? n1478 ? n1475 ? n709 ? 1'b1 : 1'b0 : 1'b0 : 1'b1 : n1478 ? n1475 ? n709 ? 1'b1 : 1'b0 : 1'b0 : n709 ? 1'b0 : 1'b1;
assign n3044 = /* LUT   22 21  6 */ n140 ? 1'b1 : 1'b0;
assign n3045 = /* LUT    5 17  3 */ n88 ? n47 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n47 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n1648 = /* LUT   21 14  0 */ n1559 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1180 ? n1632 ? 1'b0 : 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1180 ? n1632 ? 1'b0 : 1'b1 : 1'b1;
assign n3047 = /* LUT   20 26  2 */ n158 ? 1'b1 : 1'b0;
assign n3048 = /* LUT   14 20  7 */ n868 ? n526 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n526 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n751  = /* LUT   14  9  4 */ n657 ? n750 ? 1'b1 : n151 ? 1'b1 : 1'b0 : n750 ? n151 ? 1'b0 : 1'b1 : 1'b0;
assign n3050 = /* LUT   17 20  0 */ n398 ? 1'b0 : 1'b1;
assign n1487 = /* LUT   19 18  1 */ n1341 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1291 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1291 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3052 = /* LUT   10 10  3 */ n289 ? 1'b1 : 1'b0;
assign n3053 = /* LUT   23 15  7 */ n218 ? 1'b1 : 1'b0;
assign n1664 = /* LUT   21 16  3 */ n1583 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1429 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1429 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3055 = /* LUT   15 10  6 */ n763 ? 1'b1 : 1'b0;
assign n3056 = /* LUT   18 22  3 */ n272 ? n1399 ? 1'b0 : n697 ? n1273 ? 1'b0 : 1'b1 : 1'b0 : n1399 ? 1'b1 : n697 ? n1273 ? 1'b0 : 1'b1 : 1'b0;
assign n3057 = /* LUT   11 19  3 */ n260 ? 1'b0 : 1'b1;
assign n3058 = /* LUT    9 12  7 */ n155 ? n75 ? n80 ? 1'b0 : 1'b1 : 1'b1 : n75 ? n80 ? 1'b0 : 1'b1 : 1'b0;
assign n3059 = /* LUT   22 15  3 */ n59 ? 1'b0 : n802 ? n244 ? 1'b0 : n238 ? 1'b1 : 1'b0 : 1'b0;
assign n3060 = /* LUT   13 17  1 */ n494 ? 1'b0 : n184 ? 1'b0 : n345 ? 1'b0 : n185 ? 1'b0 : 1'b1;
assign n3061 = /* LUT   15 23  0 */ n1013 ? 1'b1 : 1'b0;
assign n3062 = /* LUT   18 21  7 */ n883 ? n1127 ? n46 ? 1'b1 : n731 ? 1'b0 : 1'b1 : 1'b1 : n1127 ? n46 ? n731 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n1452 = /* LUT   19 14  4 */ n967 ? n1451 ? n575 ? 1'b1 : 1'b0 : n790 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1451 ? 1'b0 : n790 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n3064 = /* LUT   22 20  5 */ n44 ? 1'b1 : 1'b0;
assign n3065 = /* LUT    5 18  2 */ n95 ? n54 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n54 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3066 = /* LUT   16 24  6 */ n32 ? 1'b1 : 1'b0;
assign n3067 = /* LUT   10 20  6 */ n159 ? 1'b1 : 1'b0;
assign n3068 = /* LUT   20 25  3 */ n42 ? 1'b1 : 1'b0;
assign n3069 = /* LUT   20 12  7 */ n218 ? 1'b1 : 1'b0;
assign n3070 = /* LUT   19 19  2 */ n42 ? 1'b1 : 1'b0;
assign n3071 = /* LUT   10 13  2 */ n307 ? n207 ? 1'b0 : n120 ? 1'b0 : 1'b1 : n207 ? n120 ? 1'b0 : 1'b1 : 1'b0;
assign n3072 = /* LUT   23 12  6 */ n140 ? 1'b1 : 1'b0;
assign n3073 = /* LUT    7 10  3 */ n111 ? n109 ? n108 ? 1'b0 : 1'b1 : 1'b1 : n109 ? 1'b0 : n108 ? 1'b1 : 1'b0;
assign n3074 = /* LUT   21 17  0 */ n1585 ? n1484 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1484 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3075 = /* LUT   15 11  5 */ n920 ? 1'b1 : 1'b0;
assign n3076 = /* LUT   18 25  2 */ n1418 ? n1151 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1151 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3077 = /* LUT   17  7  0 */ 1'b0 ? 1'b1 : 1'b0;
assign n3078 = /* LUT   20 15  3 */ n238 ? n244 ? 1'b0 : n180 ? 1'b0 : n1302 ? 1'b1 : 1'b0 : 1'b0;
assign n3079 = /* LUT   17 10  7 */ 1'b0 ? 1'b1 : 1'b0;
assign n3080 = /* LUT   22 14  4 */ n35 ? 1'b1 : 1'b0;
assign n3081 = /* LUT   13 18  0 */ n385 ? 1'b0 : 1'b1;
assign n3083 = /* LUT   15 20  1 */ n837 ? 1'b0 : 1'b1;
assign n3084 = /* LUT   18 20  4 */ n1250 ? n1383 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1383 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3085 = /* LUT   11 14  1 */ n451 ? n432 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n432 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n3086 = /* LUT   16  7  2 */ n1049 ? n902 ? 1'b0 : n737 ? 1'b0 : 1'b1 : n902 ? n737 ? 1'b0 : 1'b1 : 1'b0;
assign n3087 = /* LUT   19 15  7 */ n1322 ? n1465 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1465 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3088 = /* LUT   22 23  4 */ n35 ? 1'b1 : 1'b0;
assign n3089 = /* LUT   15 26  0 */ n1043 ? n898 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n898 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3090 = /* LUT   12 12  2 */ n426 ? 1'b1 : 1'b0;
assign n3091 = /* LUT   17 22  2 */ n980 ? 1'b0 : 1'b1;
assign n3092 = /* LUT   14 11  6 */ n662 ? 1'b1 : 1'b0;
assign n3093 = /* LUT   19 16  3 */ n42 ? 1'b1 : 1'b0;
assign n3094 = /* LUT   10 12  1 */ n43 ? n136 ? 1'b0 : n196 ? 1'b1 : 1'b0 : 1'b1;
assign n3095 = /* LUT   22 10  1 */ n1701 ? n1622 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n1622 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3096 = /* LUT   21 18  1 */ n1366 ? n1673 ? n575 ? 1'b1 : 1'b0 : n810 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1673 ? 1'b0 : n810 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n3097 = /* LUT   12 15  4 */ n499 ? 1'b0 : 1'b1;
assign n3098 = /* LUT   18 24  1 */ n1035 ? n575 ? n644 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n644 ? 1'b1 : 1'b0 : 1'b0;
assign n908  = /* LUT   15  7  5 */ n651 ? 1'b0 : n646 ? n649 ? 1'b0 : n650 ? 1'b0 : 1'b1 : 1'b0;
assign n1567 = /* LUT   20 14  0 */ n1447 ? n709 ? n1560 ? 1'b1 : 1'b0 : 1'b0 : n709 ? n1105 ? 1'b1 : 1'b0 : 1'b1;
assign n3100 = /* LUT   13  8  6 */ n149 ? n653 ? 1'b1 : n648 ? 1'b1 : 1'b0 : n653 ? n648 ? 1'b0 : 1'b1 : 1'b0;
assign n3101 = /* LUT   13 19  7 */ n513 ? 1'b0 : 1'b1;
assign n3102 = /* LUT   18 23  5 */ n47 ? n1127 ? n887 ? 1'b1 : n731 ? 1'b1 : 1'b0 : n887 ? 1'b1 : 1'b0 : n1127 ? n887 ? n731 ? 1'b0 : 1'b1 : 1'b0 : n887 ? 1'b1 : 1'b0;
assign n3103 = /* LUT   14 18  6 */ n833 ? n185 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n185 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n3104 = /* LUT   11 15  2 */ n475 ? n297 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n297 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n3105 = /* LUT   14  7  1 */ n741 ? n647 ? 1'b0 : n734 ? 1'b0 : 1'b1 : n647 ? n734 ? 1'b0 : 1'b1 : 1'b0;
assign n1435 = /* LUT   19 12  6 */ n59 ? n440 ? 1'b1 : 1'b0 : 1'b0;
assign n3106 = /* LUT   12 19  3 */ n42 ? 1'b1 : 1'b0;
assign n3107 = /* LUT   14 17  0 */ n398 ? 1'b0 : n526 ? 1'b0 : n528 ? 1'b0 : n527 ? 1'b0 : 1'b1;
assign n3108 = /* LUT   17 12  4 */ n940 ? n928 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n928 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3109 = /* LUT   17 23  5 */ n988 ? 1'b0 : 1'b1;
assign n3110 = /* LUT   10 15  0 */ io_0_25_1 ? n214 ? 1'b1 : 1'b0 : 1'b0;
assign n3112 = /* LUT   21 19  6 */ n712 ? n1684 ? 1'b1 : 1'b0 : n1608 ? 1'b1 : 1'b0;
assign n3115 = /* LUT   15  9  3 */ n735 ? 1'b1 : 1'b0;
assign n3116 = /* LUT   12 14  7 */ n491 ? 1'b0 : 1'b1;
assign n3117 = /* LUT    6 16  0 */ io_0_20_0 ? 1'b0 : io_0_16_0 ? 1'b0 : io_25_0_0 ? 1'b0 : 1'b1;
assign n1557 = /* LUT   20 13  1 */ n1439 ? n1541 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1541 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3119 = /* LUT   16 23  1 */ io_8_33_0 ? 1'b1 : 1'b0;
assign n3120 = /* LUT   10 17  4 */ n363 ? n227 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n227 ? 1'b1 : 1'b0;
assign n3121 = /* LUT   13 20  6 */ n190 ? 1'b0 : 1'b1;
assign n1314 = /* LUT   18 13  3 */ n1084 ? n1313 ? n709 ? 1'b1 : 1'b0 : n1310 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1313 ? 1'b0 : n1310 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n3123 = /* LUT   20 19  0 */ n159 ? 1'b1 : 1'b0;
assign n3124 = /* LUT   14 13  7 */ n218 ? 1'b1 : 1'b0;
assign n3125 = /* LUT   11 12  3 */ n427 ? 1'b1 : 1'b0;
assign n1443 = /* LUT   19 13  1 */ n1427 ? n1180 ? 1'b0 : n575 ? 1'b1 : n1422 ? 1'b0 : 1'b1 : n1180 ? n575 ? 1'b0 : 1'b1 : n575 ? 1'b1 : n1422 ? 1'b0 : 1'b1;
assign n1731 = /* LUT   22 17  2 */ n1492 ? n709 ? n930 ? 1'b0 : 1'b1 : n1473 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1473 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n3130 = /* LUT   15 24  2 */ n1028 ? n884 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n884 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3131 = /* LUT   12 18  0 */ n604 ? n484 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n484 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3132 = /* LUT   17 13  7 */ n450 ? n1189 ? 1'b1 : n575 ? 1'b1 : 1'b0 : n1189 ? n575 ? 1'b0 : 1'b1 : 1'b0;
assign n3133 = /* LUT   14 16  3 */ n696 ? 1'b1 : 1'b0;
assign n1213 = /* LUT   17 16  4 */ n1075 ? n575 ? n1164 ? 1'b1 : 1'b0 : 1'b0 : n575 ? n1211 ? 1'b1 : 1'b0 : 1'b1;
assign n3135 = /* LUT    7  9  6 */ n64 ? 1'b1 : n108 ? n109 ? 1'b0 : 1'b1 : n65 ? 1'b1 : 1'b0;
assign n3136 = /* LUT   21 20  7 */ n218 ? 1'b1 : 1'b0;
assign n3139 = /* LUT   15 14  2 */ n244 ? 1'b0 : n956 ? 1'b1 : 1'b0;
assign n3140 = /* LUT   18 17  6 */ n1350 ? n1354 ? n709 ? 1'b1 : 1'b0 : n1230 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1354 ? 1'b0 : n1230 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n3141 = /* LUT   12 13  6 */ n140 ? 1'b1 : 1'b0;
assign n3142 = /* LUT   16 22  2 */ n1127 ? n892 ? n53 ? 1'b1 : n731 ? 1'b0 : 1'b1 : n53 ? n731 ? 1'b1 : 1'b0 : 1'b0 : n892 ? 1'b1 : 1'b0;
assign n3143 = /* LUT   10 16  7 */ n352 ? n237 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n237 ? 1'b1 : 1'b0;
assign n3144 = /* LUT   13 10  4 */ n669 ? 1'b1 : 1'b0;
assign n3145 = /* LUT   18 12  0 */ n159 ? 1'b1 : 1'b0;
assign n773  = /* LUT   14 12  4 */ n770 ? 1'b0 : io_0_25_1 ? n771 ? n591 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3147 = /* LUT   11 13  4 */ n140 ? 1'b1 : 1'b0;
assign n3148 = /* LUT   19 10  0 */ n159 ? 1'b1 : 1'b0;
assign n1722 = /* LUT   22 16  1 */ n1647 ? n575 ? n1180 ? 1'b0 : 1'b1 : n574 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n574 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3150 = /* LUT   15 25  5 */ n1040 ? n885 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n885 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3151 = /* LUT   12 17  1 */ n597 ? n469 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n469 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3152 = /* LUT   14 19  2 */ n846 ? n516 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n516 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n1198 = /* LUT   17 14  6 */ n1096 ? n575 ? n1180 ? 1'b0 : 1'b1 : n695 ? 1'b0 : n1180 ? 1'b0 : 1'b1 : n575 ? n1180 ? 1'b0 : 1'b1 : n695 ? n1180 ? 1'b1 : 1'b0 : 1'b1;
assign n3154 = /* LUT   17 17  7 */ n709 ? n595 ? 1'b1 : 1'b0 : n930 ? n595 ? n575 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3155 = /* LUT   21 21  4 */ n1690 ? n575 ? n1691 ? 1'b1 : 1'b0 : 1'b1 : n575 ? n1691 ? 1'b1 : 1'b0 : 1'b0;
assign n3156 = /* LUT   15 15  1 */ n212 ? 1'b1 : 1'b0;
assign n3157 = /* LUT   11  9  1 */ n280 ? 1'b0 : n406 ? n281 ? 1'b0 : 1'b1 : 1'b0;
assign n3158 = /* LUT   16 21  3 */ n158 ? 1'b1 : 1'b0;
assign n3159 = /* LUT   10 19  6 */ n140 ? 1'b1 : 1'b0;
assign n3160 = /* LUT   13 11  3 */ n565 ? io_33_1_1 ? n560 ? 1'b0 : 1'b1 : n561 ? 1'b0 : n560 ? 1'b0 : 1'b1 : io_33_1_1 ? n560 ? 1'b1 : 1'b0 : n561 ? 1'b0 : n560 ? 1'b1 : 1'b0;
assign n3161 = /* LUT   13 22  4 */ n402 ? 1'b0 : 1'b1;
assign n3162 = /* LUT   18 15  1 */ n159 ? 1'b1 : 1'b0;
assign n3163 = /* LUT   20 17  2 */ n1470 ? n1483 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1483 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n798  = /* LUT   14 15  5 */ n696 ? n578 ? 1'b0 : n577 ? n579 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3164 = /* LUT   11 10  5 */ n65 ? 1'b0 : n194 ? n411 ? 1'b1 : 1'b0 : n409 ? 1'b1 : 1'b0;
assign n3165 = /* LUT   19 11  3 */ n42 ? 1'b1 : 1'b0;
assign n3166 = /* LUT   17 15  1 */ n1103 ? n1205 ? n575 ? 1'b1 : 1'b0 : n1203 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1205 ? 1'b0 : n1203 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n3167 = /* LUT   19 25  0 */ n159 ? 1'b1 : 1'b0;
assign n3170 = /* LUT   22 13  4 */ n1308 ? n1714 ? n575 ? 1'b1 : 1'b0 : n1549 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1714 ? 1'b0 : n1549 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n3171 = /* LUT   21 22  5 */ n1604 ? n1698 ? 1'b1 : n575 ? 1'b1 : 1'b0 : n1698 ? n575 ? 1'b0 : 1'b1 : 1'b0;
assign n3172 = /* LUT   15 12  0 */ n769 ? n126 ? n159 ? 1'b1 : n592 ? 1'b0 : 1'b1 : n159 ? n592 ? 1'b1 : 1'b0 : 1'b0 : n126 ? 1'b1 : 1'b0;
assign n3173 = /* LUT   18 19  4 */ n1373 ? n823 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n823 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3174 = /* LUT   11 22  0 */ n159 ? 1'b1 : 1'b0;
assign n3175 = /* LUT   16 15  5 */ n948 ? n244 ? n525 ? 1'b0 : n59 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n3176 = /* LUT   16 20  4 */ n59 ? n936 ? n540 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3177 = /* LUT   13 12  2 */ n679 ? 1'b1 : 1'b0;
assign n3178 = /* LUT   15 18  3 */ n42 ? 1'b1 : 1'b0;
assign n3179 = /* LUT   20 16  5 */ n158 ? 1'b1 : 1'b0;
assign n3180 = /* LUT   12 20  3 */ n42 ? 1'b1 : 1'b0;
assign n3181 = /* LUT   17 11  6 */ n158 ? 1'b1 : 1'b0;
assign n3182 = /* LUT   11 11  6 */ n421 ? n295 ? 1'b0 : n282 ? 1'b0 : 1'b1 : n295 ? n282 ? 1'b0 : 1'b1 : 1'b0;
assign n3183 = /* LUT   23 14  3 */ n42 ? 1'b1 : 1'b0;
assign n1628 = /* LUT   21 10  0 */ n1536 ? n1535 ? 1'b0 : n1624 ? 1'b0 : 1'b1 : 1'b0;
assign n3186 = /* LUT   19 22  1 */ n1511 ? n1390 ? 1'b0 : n1258 ? 1'b0 : 1'b1 : n1390 ? n1258 ? 1'b0 : 1'b1 : 1'b0;
assign n3187 = /* LUT   16 16  1 */ n212 ? 1'b1 : 1'b0;
assign n3188 = /* LUT   22 12  7 */ n218 ? 1'b1 : 1'b0;
assign n3189 = /* LUT    7 12  5 */ n43 ? 1'b0 : 1'b1;
assign n3190 = /* LUT   18 18  3 */ n158 ? 1'b1 : 1'b0;
assign n3191 = /* LUT   20 20  2 */ n44 ? 1'b1 : 1'b0;
assign n3192 = /* LUT   14 10  7 */ n759 ? 1'b1 : 1'b0;
assign n3193 = /* LUT   16 14  6 */ n59 ? 1'b0 : n1086 ? n244 ? 1'b0 : n525 ? 1'b0 : 1'b1 : 1'b0;
assign n3194 = /* LUT    5 17  4 */ n89 ? n48 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n48 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3195 = /* LUT   16 19  5 */ n218 ? 1'b1 : 1'b0;
assign n3196 = /* LUT   15 19  0 */ n159 ? 1'b1 : 1'b0;
assign n750  = /* LUT   14  9  3 */ n152 ? n749 ? 1'b1 : 1'b0 : n665 ? 1'b1 : 1'b0;
assign n3198 = /* LUT   17 20  7 */ n526 ? 1'b0 : 1'b1;
assign n3199 = /* LUT   23 15  0 */ n159 ? 1'b1 : 1'b0;
assign n3200 = /* LUT   24 16  0 */ n44 ? 1'b1 : 1'b0;
assign n1666 = /* LUT   21 16  6 */ n685 ? n1665 ? 1'b1 : n575 ? 1'b1 : 1'b0 : n1665 ? n575 ? 1'b0 : 1'b1 : 1'b0;
assign n3202 = /* LUT   21 11  7 */ n218 ? 1'b1 : 1'b0;
assign n3205 = /* LUT   19 23  2 */ n1025 ? io_0_25_1 ? n272 ? n729 ? 1'b1 : 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n3206 = /* LUT   22 15  6 */ n238 ? n244 ? 1'b0 : n525 ? 1'b0 : n59 ? 1'b0 : 1'b1 : 1'b0;
assign n3207 = /* LUT   18 21  2 */ n882 ? n30 ? 1'b1 : n731 ? n1127 ? 1'b0 : 1'b1 : 1'b1 : n30 ? n731 ? n1127 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3208 = /* LUT   20 11  3 */ n35 ? 1'b1 : 1'b0;
assign n3209 = /* LUT   11 20  2 */ n249 ? 1'b0 : 1'b1;
assign n3210 = /* LUT   16 13  7 */ n244 ? n1079 ? 1'b0 : n590 ? 1'b1 : 1'b0 : 1'b0;
assign n3211 = /* LUT    5 18  5 */ n98 ? n57 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n57 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3212 = /* LUT   16 18  6 */ n140 ? 1'b1 : 1'b0;
assign n3213 = /* LUT   10 20  3 */ n158 ? 1'b1 : 1'b0;
assign n3214 = /* LUT   15 16  1 */ n238 ? n244 ? 1'b0 : n59 ? n525 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n3215 = /* LUT   21 15  4 */ n1575 ? n1658 ? n930 ? 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? 1'b0 : 1'b1 : n1658 ? n930 ? n709 ? 1'b1 : 1'b0 : n709 ? 1'b0 : 1'b1 : n930 ? n709 ? 1'b1 : 1'b0 : 1'b1;
assign n3216 = /* LUT   20 25  6 */ n140 ? 1'b1 : 1'b0;
assign n3217 = /* LUT   20 22  7 */ io_11_33_1 ? n994 ? 1'b1 : 1'b0 : 1'b1;
assign n3220 = /* LUT   23 12  1 */ n212 ? 1'b1 : 1'b0;
assign n3221 = /* LUT   24 15  1 */ n212 ? 1'b1 : 1'b0;
assign n3222 = /* LUT    7 10  6 */ n41 ? 1'b1 : 1'b0;
assign n3223 = /* LUT   21 17  5 */ n158 ? 1'b1 : 1'b0;
assign n3224 = /* LUT   21 12  6 */ n140 ? 1'b1 : 1'b0;
assign n3225 = /* LUT   12 21  5 */ n521 ? 1'b0 : 1'b1;
assign n3226 = /* LUT   17 10  2 */ 1'b0 ? 1'b1 : 1'b0;
assign n3227 = /* LUT   19 20  3 */ n272 ? n1379 ? io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0;
assign n3228 = /* LUT   22 14  1 */ n212 ? 1'b1 : 1'b0;
assign n1386 = /* LUT   18 20  1 */ n1280 ? n1385 ? n709 ? n930 ? 1'b0 : 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n1385 ? n709 ? n930 ? 1'b0 : 1'b1 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n3230 = /* LUT   20 10  0 */ n1539 ? n41 ? n1540 ? 1'b1 : 1'b0 : n1537 ? n1540 ? 1'b1 : 1'b0 : 1'b0 : n41 ? 1'b1 : n1537 ? n1540 ? 1'b1 : 1'b0 : 1'b0;
assign n3231 = /* LUT   23 16  7 */ n218 ? 1'b1 : 1'b0;
assign n3232 = /* LUT   11 14  4 */ n454 ? n435 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n435 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n3233 = /* LUT   16 12  0 */ n440 ? 1'b1 : n180 ? 1'b1 : 1'b0;
assign n3234 = /* LUT    5 19  2 */ n103 ? n30 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n30 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3235 = /* LUT   16 17  7 */ n218 ? 1'b1 : 1'b0;
assign n3236 = /* LUT   15 17  6 */ n140 ? 1'b1 : 1'b0;
assign n3237 = /* LUT   20 24  1 */ n1519 ? n1406 ? n1405 ? n1518 ? 1'b1 : 1'b0 : n1518 ? 1'b0 : 1'b1 : 1'b0 : n1406 ? 1'b0 : n1405 ? n1518 ? 1'b1 : 1'b0 : n1518 ? 1'b0 : 1'b1;
assign n3238 = /* LUT   12 12  7 */ n424 ? 1'b1 : 1'b0;
assign n3239 = /* LUT   20 21  6 */ n1499 ? n1505 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1505 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3240 = /* LUT   17 22  5 */ n844 ? 1'b0 : 1'b1;
assign n3241 = /* LUT   24 14  2 */ n44 ? 1'b1 : 1'b0;
assign n3242 = /* LUT   22 10  6 */ n1706 ? n1626 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n1626 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3243 = /* LUT   21 18  4 */ n1367 ? n1674 ? n575 ? 1'b1 : 1'b0 : n811 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1674 ? 1'b0 : n811 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n1645 = /* LUT   21 13  5 */ n1563 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1428 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1428 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3245 = /* LUT   12 15  3 */ n487 ? 1'b0 : 1'b1;
assign n3246 = /* LUT   19 21  4 */ n1025 ? 1'b0 : n1242 ? n641 ? 1'b1 : n1388 ? 1'b1 : 1'b0 : n641 ? 1'b0 : n1388 ? 1'b1 : 1'b0;
assign n3247 = /* LUT   10 11  0 */ n291 ? n201 ? 1'b0 : 1'b1 : n201 ? 1'b1 : 1'b0;
assign n3248 = /* LUT   15 21  3 */ n999 ? 1'b0 : 1'b1;
assign n3249 = /* LUT   18 23  0 */ n731 ? n886 ? n1127 ? n45 ? 1'b1 : 1'b0 : 1'b1 : n1127 ? n45 ? 1'b1 : 1'b0 : 1'b0 : n886 ? 1'b1 : 1'b0;
assign n3250 = /* LUT   23 17  0 */ n42 ? 1'b1 : 1'b0;
assign n3251 = /* LUT   11 15  7 */ n480 ? n302 ? 1'b1 : 1'b0 : n302 ? 1'b0 : 1'b1;
assign n3252 = /* LUT   14  7  4 */ n744 ? n650 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n650 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3253 = /* LUT   11 18  4 */ n507 ? 1'b0 : 1'b1;
assign n3254 = /* LUT   16 11  1 */ n212 ? 1'b1 : 1'b0;
assign n3257 = /* LUT   18  9  3 */ n1284 ? 1'b1 : 1'b0;
assign n3258 = /* LUT   12 19  6 */ n140 ? 1'b1 : 1'b0;
assign n3259 = /* LUT    6 11  6 */ n118 ? n73 ? 1'b0 : n81 ? 1'b0 : 1'b1 : n73 ? n81 ? 1'b0 : 1'b1 : 1'b0;
assign n3260 = /* LUT   17 23  2 */ n878 ? 1'b0 : 1'b1;
assign n1477 = /* LUT   19 17  1 */ n1347 ? n1476 ? n705 ? 1'b0 : 1'b1 : 1'b0 : n1357 ? 1'b1 : n705 ? 1'b1 : 1'b0;
assign n3262 = /* LUT   22 21  2 */ n44 ? 1'b1 : 1'b0;
assign n1682 = /* LUT   21 19  3 */ n1330 ? n709 ? n930 ? 1'b0 : 1'b1 : n1580 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1580 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n3264 = /* LUT   21 14  4 */ n1432 ? n1649 ? n575 ? 1'b1 : 1'b0 : n1546 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1649 ? 1'b0 : n1546 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n3265 = /* LUT    9 16  1 */ n241 ? n242 ? n243 ? n240 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n3266 = /* LUT   12 14  0 */ n468 ? 1'b0 : 1'b1;
assign n3268 = /* LUT   14 20  3 */ n864 ? n527 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n527 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n3269 = /* LUT   19 18  5 */ n1358 ? n1489 ? n1058 ? n709 ? 1'b0 : 1'b1 : 1'b1 : n1058 ? 1'b0 : 1'b1 : n1489 ? n1058 ? n709 ? 1'b0 : 1'b1 : n709 ? 1'b1 : 1'b0 : n1058 ? 1'b0 : n709 ? 1'b1 : 1'b0;
assign n3272 = /* LUT   16 23  4 */ io_0_11_1 ? 1'b1 : 1'b0;
assign n3273 = /* LUT   15 10  2 */ n766 ? 1'b1 : 1'b0;
assign n3274 = /* LUT   20 19  7 */ n218 ? 1'b1 : 1'b0;
assign n3275 = /* LUT   20  8  6 */ 1'b0 ? 1'b1 : 1'b0;
assign n3276 = /* LUT   11 12  6 */ n423 ? 1'b1 : 1'b0;
assign n3279 = /* LUT   11 19  7 */ n264 ? 1'b0 : 1'b1;
assign n3280 = /* LUT   16 10  2 */ n1055 ? 1'b1 : 1'b0;
assign n3281 = /* LUT    9 12  3 */ n155 ? 1'b1 : n205 ? 1'b0 : n43 ? 1'b1 : 1'b0;
assign n3282 = /* LUT   15 24  5 */ n1031 ? n889 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n889 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3283 = /* LUT   12 18  5 */ n614 ? n488 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n488 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3284 = /* LUT   17 16  3 */ n1194 ? n1212 ? n575 ? n1193 ? 1'b1 : 1'b0 : 1'b0 : 1'b1 : n1212 ? n575 ? n1193 ? 1'b1 : 1'b0 : 1'b0 : n575 ? 1'b0 : 1'b1;
assign n3285 = /* LUT   19 14  0 */ n158 ? 1'b1 : 1'b0;
assign n3286 = /* LUT   22 20  1 */ n1686 ? n1692 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1692 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3287 = /* LUT   16 24  2 */ io_6_33_0 ? 1'b1 : 1'b0;
assign n3288 = /* LUT   21 20  2 */ n44 ? 1'b1 : 1'b0;
assign n3289 = /* LUT   12 13  1 */ n212 ? 1'b1 : 1'b0;
assign n3290 = /* LUT   14 23  2 */ n35 ? 1'b1 : 1'b0;
assign n3291 = /* LUT   20 12  3 */ n42 ? 1'b1 : 1'b0;
assign n3292 = /* LUT   19 19  6 */ n218 ? 1'b1 : 1'b0;
assign n3293 = /* LUT   10 13  6 */ n311 ? n210 ? 1'b0 : n120 ? 1'b0 : 1'b1 : n210 ? n120 ? 1'b0 : 1'b1 : 1'b0;
assign n3294 = /* LUT   15 11  1 */ n660 ? 1'b1 : 1'b0;
assign n3295 = /* LUT   20 18  4 */ n212 ? 1'b1 : 1'b0;
assign n3296 = /* LUT   20 15  7 */ n592 ? n590 ? n244 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3297 = /* LUT   11 13  1 */ n42 ? 1'b1 : 1'b0;
assign n3298 = /* LUT   11 16  6 */ n358 ? 1'b1 : 1'b0;
assign n3299 = /* LUT   13  7  3 */ io_33_1_1 ? 1'b0 : n656 ? n544 ? 1'b1 : n646 ? 1'b0 : 1'b1 : n544 ? n646 ? 1'b1 : 1'b0 : 1'b0;
assign n3300 = /* LUT   15 25  2 */ n1037 ? n894 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n894 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3301 = /* LUT   18 11  1 */ n212 ? 1'b1 : 1'b0;
assign n3302 = /* LUT   15 20  5 */ n840 ? 1'b0 : 1'b1;
assign n3303 = /* LUT   12 17  4 */ n600 ? n472 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n472 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3304 = /* LUT   17 17  0 */ n1091 ? n575 ? n1108 ? 1'b1 : 1'b0 : 1'b0 : n575 ? n809 ? 1'b1 : 1'b0 : 1'b1;
assign n1464 = /* LUT   19 15  3 */ n1340 ? n1462 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1462 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n3306 = /* LUT   22 23  0 */ n159 ? 1'b1 : 1'b0;
assign n1696 = /* LUT   21 21  1 */ n1279 ? n1695 ? n709 ? n930 ? 1'b0 : 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n1695 ? n709 ? n930 ? 1'b0 : 1'b1 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n3308 = /* LUT    9 18  3 */ n218 ? 1'b1 : 1'b0;
assign n3309 = /* LUT   14 22  5 */ n218 ? 1'b1 : 1'b0;
assign n408  = /* LUT   11  9  6 */ n152 ? n276 ? n151 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3310 = /* LUT   19 16  7 */ n218 ? 1'b1 : 1'b0;
assign n3311 = /* LUT   16 21  6 */ n159 ? 1'b1 : 1'b0;
assign n912  = /* LUT   15  8  0 */ n746 ? n911 ? 1'b1 : n648 ? 1'b1 : 1'b0 : n911 ? n648 ? 1'b0 : 1'b1 : 1'b0;
assign n3313 = /* LUT   20 17  5 */ n44 ? 1'b1 : 1'b0;
assign n123  = /* LUT    6 12  4 */ n72 ? 1'b1 : n74 ? 1'b1 : n73 ? 1'b1 : n71 ? 1'b1 : 1'b0;
assign n1570 = /* LUT   20 14  4 */ n1068 ? n1569 ? n709 ? 1'b1 : 1'b0 : n1564 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1569 ? 1'b0 : n1564 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n3315 = /* LUT   23 20  3 */ n42 ? 1'b1 : 1'b0;
assign n412  = /* LUT   11 10  0 */ n284 ? n154 ? 1'b0 : 1'b1 : 1'b1;
assign n3316 = /* LUT   14 18  2 */ n829 ? n386 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n386 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n3319 = /* LUT   19 12  2 */ n802 ? n244 ? 1'b0 : n59 ? 1'b0 : n590 ? 1'b1 : 1'b0 : 1'b0;
assign n3320 = /* LUT   21 22  0 */ n1700 ? n1533 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1533 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3321 = /* LUT   17 12  0 */ n140 ? 1'b1 : 1'b0;
assign n818  = /* LUT   14 17  4 */ n713 ? n817 ? n705 ? 1'b0 : 1'b1 : n794 ? 1'b1 : n705 ? 1'b1 : 1'b0 : n817 ? 1'b0 : n794 ? 1'b1 : n705 ? 1'b1 : 1'b0;
assign n3323 = /* LUT   11 22  7 */ n42 ? 1'b1 : 1'b0;
assign n3324 = /* LUT   10 15  4 */ n335 ? n223 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n223 ? 1'b1 : 1'b0;
assign n3325 = /* LUT   16 20  1 */ n238 ? n157 ? n244 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3326 = /* LUT   15 18  6 */ n140 ? 1'b1 : 1'b0;
assign n3329 = /* LUT   18 14  3 */ n1092 ? n1325 ? n709 ? 1'b1 : 1'b0 : n1090 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1325 ? 1'b0 : n1090 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n3330 = /* LUT   20 16  2 */ n44 ? 1'b1 : 1'b0;
assign n3331 = /* LUT   20 13  5 */ n212 ? 1'b1 : 1'b0;
assign n3332 = /* LUT   11 11  3 */ n418 ? n286 ? 1'b0 : n282 ? 1'b0 : 1'b1 : n286 ? n282 ? 1'b0 : 1'b1 : 1'b0;
assign n1738 = /* LUT   22 18  4 */ n1495 ? n709 ? n930 ? 1'b0 : 1'b1 : n1735 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n1735 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n3334 = /* LUT   10 17  0 */ n353 ? n242 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n242 ? 1'b1 : 1'b0;
assign n3335 = /* LUT    9 15  6 */ n170 ? n230 ? n44 ? 1'b0 : n35 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n3336 = /* LUT   18 13  7 */ n1087 ? n1315 ? n709 ? 1'b1 : 1'b0 : n1081 ? 1'b1 : n709 ? 1'b0 : 1'b1 : n1315 ? 1'b0 : n1081 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n3339 = /* LUT   14 13  3 */ n42 ? 1'b1 : 1'b0;
assign n3340 = /* LUT   19 22  4 */ n1514 ? n1393 ? 1'b0 : n1258 ? 1'b0 : 1'b1 : n1393 ? n1258 ? 1'b0 : 1'b1 : 1'b0;
assign n1445 = /* LUT   19 13  5 */ n1434 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1289 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1289 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3342 = /* LUT   22 17  6 */ n1667 ? n705 ? n595 ? n1672 ? 1'b0 : 1'b1 : 1'b0 : n595 ? 1'b0 : 1'b1 : n705 ? n595 ? n1672 ? 1'b0 : 1'b1 : 1'b1 : n595 ? 1'b0 : 1'b1;
assign n3343 = /* LUT   16 16  6 */ n140 ? 1'b1 : 1'b0;
assign n947  = /* LUT   15 13  4 */ n778 ? 1'b1 : n689 ? n943 ? n779 ? 1'b0 : 1'b1 : 1'b1 : 1'b1;
assign n3344 = /* LUT   20 20  7 */ n218 ? 1'b1 : 1'b0;
assign n3345 = /* LUT   14 16  7 */ n547 ? 1'b1 : 1'b0;
assign n1188 = /* LUT   17 13  3 */ n1065 ? n709 ? n1066 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n709 ? n1066 ? n930 ? 1'b0 : 1'b1 : 1'b1 : n930 ? 1'b0 : 1'b1;
assign n3347 = /* LUT   16 19  0 */ n44 ? 1'b1 : 1'b0;
assign n3348 = /* LUT    9 11  3 */ n7 ? 1'b1 : io_0_25_1 ? 1'b1 : 1'b0;
assign n3349 = /* LUT   15 19  5 */ n158 ? 1'b1 : 1'b0;
assign n3352 = /* LUT   18 17  2 */ n1241 ? n1352 ? n709 ? 1'b1 : 1'b0 : 1'b0 : n1215 ? 1'b1 : n709 ? 1'b0 : 1'b1;
assign n957  = /* LUT   15 14  6 */ n771 ? 1'b0 : n770 ? 1'b1 : 1'b0;
assign n3353 = /* LUT   20 23  3 */ n212 ? 1'b1 : 1'b0;
assign n3354 = /* LUT   10 16  3 */ n348 ? n233 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n233 ? 1'b1 : 1'b0;
assign n3355 = /* LUT   13 10  0 */ n668 ? 1'b1 : 1'b0;
assign n3356 = /* LUT   18 12  4 */ n35 ? 1'b1 : 1'b0;
assign n772  = /* LUT   14 12  0 */ n671 ? n152 ? n670 ? 1'b1 : 1'b0 : 1'b1 : n152 ? n670 ? 1'b1 : 1'b0 : 1'b0;
assign n3360 = /* LUT   19 23  7 */ n272 ? n1148 ? io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : io_0_25_1 ? n1025 ? 1'b1 : 1'b0 : 1'b0;
assign n3361 = /* LUT   19 10  4 */ n35 ? 1'b1 : 1'b0;
assign n1724 = /* LUT   22 16  5 */ n1590 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1426 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1426 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3363 = /* LUT   20 11  6 */ n218 ? 1'b1 : 1'b0;
assign n3364 = /* LUT   17 14  2 */ n158 ? 1'b1 : 1'b0;
assign n3365 = /* LUT   14 19  6 */ n850 ? n188 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n188 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n3366 = /* LUT   19 24  3 */ n1528 ? n1408 ? 1'b0 : n1501 ? 1'b0 : 1'b1 : n1408 ? n1501 ? 1'b0 : 1'b1 : 1'b0;
assign n3367 = /* LUT   11 20  5 */ n252 ? 1'b0 : 1'b1;
assign n3368 = /* LUT   16 18  3 */ n42 ? 1'b1 : 1'b0;
assign n3369 = /* LUT   15 16  4 */ n59 ? n180 ? 1'b0 : n244 ? 1'b0 : n141 ? 1'b1 : 1'b0 : 1'b0;
assign n3370 = /* LUT   15 15  5 */ n158 ? 1'b1 : 1'b0;
assign n3371 = /* LUT   18 16  1 */ n1342 ? n709 ? 1'b0 : n712 ? 1'b1 : 1'b0 : n709 ? n712 ? 1'b1 : 1'b0 : 1'b0;
assign n3372 = /* LUT   20 22  0 */ n1394 ? 1'b1 : n1393 ? 1'b1 : n1396 ? 1'b1 : n1389 ? 1'b1 : 1'b0;
assign n3375 = /* LUT   10 19  2 */ n44 ? 1'b1 : 1'b0;
assign n1335 = /* LUT   18 15  5 */ n683 ? n1334 ? 1'b1 : n575 ? 1'b1 : 1'b0 : n1334 ? n575 ? 1'b0 : 1'b1 : 1'b0;
assign n3377 = /* LUT   12 21  0 */ n518 ? 1'b0 : 1'b1;
assign n3379 = /* LUT   14 15  1 */ n140 ? 1'b1 : 1'b0;
assign n3380 = /* LUT   19 20  6 */ n590 ? n157 ? n244 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3381 = /* LUT   19 11  7 */ n218 ? 1'b1 : 1'b0;
assign n3382 = /* LUT   22 19  4 */ n1677 ? n1607 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1607 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3383 = /* LUT   24 18  2 */ 1'b0 ? 1'b1 : 1'b0;
assign n1207 = /* LUT   17 15  5 */ n171 ? n575 ? n1180 ? 1'b0 : 1'b1 : n973 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n973 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3385 = /* LUT   16 17  2 */ n44 ? 1'b1 : 1'b0;
assign n1713 = /* LUT   22 13  0 */ n1639 ? n575 ? n1180 ? 1'b0 : 1'b1 : n1635 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n575 ? n1180 ? 1'b0 : 1'b1 : n1635 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3387 = /* LUT   15 17  3 */ n42 ? 1'b1 : 1'b0;
assign n3388 = /* LUT   15 12  4 */ n761 ? n152 ? n765 ? 1'b1 : 1'b0 : 1'b1 : n152 ? n765 ? 1'b1 : 1'b0 : 1'b0;
assign n3389 = /* LUT   18 19  0 */ n1233 ? n1372 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1372 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3390 = /* LUT   20 21  1 */ n42 ? 1'b1 : 1'b0;
assign n3391 = /* LUT   17 25  1 */ n712 ? n575 ? 1'b0 : 1'b1 : 1'b1;
assign n3392 = /* LUT   16 15  1 */ n244 ? 1'b0 : n1097 ? n802 ? n59 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3393 = /* LUT   23 13  3 */ n158 ? 1'b1 : 1'b0;
assign n3394 = /* LUT   24 14  7 */ n218 ? 1'b1 : 1'b0;
assign n3395 = /* LUT   17 11  2 */ n1057 ? n1168 ? n709 ? 1'b0 : n930 ? 1'b0 : 1'b1 : n930 ? 1'b0 : 1'b1 : n1168 ? n709 ? n930 ? 1'b1 : 1'b0 : n930 ? 1'b0 : 1'b1 : n709 ? 1'b1 : n930 ? 1'b0 : 1'b1;
assign n3396 = /* LUT   19 21  1 */ n641 ? n1500 ? n1025 ? 1'b0 : 1'b1 : 1'b0 : n880 ? n1025 ? 1'b0 : 1'b1 : 1'b0;
assign n3397 = /* LUT   11 17  7 */ n495 ? 1'b0 : n498 ? n179 ? n374 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3398 = /* LUT   23 14  7 */ n218 ? 1'b1 : 1'b0;
assign n3399 = /* LUT   24 17  3 */ n42 ? 1'b1 : 1'b0;
assign n3400 = /* LUT   17  8  4 */ n1158 ? 1'b1 : 1'b0;
assign n3401 = /* LUT   11 18  3 */ n506 ? 1'b0 : 1'b1;
assign n3402 = /* LUT   22 12  3 */ n42 ? 1'b1 : 1'b0;
assign n3403 = /* LUT   13 16  5 */ n218 ? 1'b1 : 1'b0;
assign n3406 = /* LUT   18  9  6 */ n1285 ? 1'b1 : 1'b0;
assign n3407 = /* LUT   18 18  7 */ n1235 ? n1365 ? n1232 ? n709 ? 1'b1 : 1'b0 : 1'b0 : 1'b1 : n1365 ? n1232 ? n709 ? 1'b1 : 1'b0 : 1'b0 : n709 ? 1'b0 : 1'b1;
assign n3408 = /* LUT    6 11  1 */ n113 ? n68 ? 1'b0 : n81 ? 1'b0 : 1'b1 : n68 ? n81 ? 1'b0 : 1'b1 : 1'b0;
assign n3409 = /* LUT   23 18  1 */ n212 ? 1'b1 : 1'b0;
assign n3410 = /* LUT   14 10  3 */ n760 ? 1'b1 : 1'b0;
assign n3411 = /* LUT   19 17  6 */ n1223 ? n1479 ? n705 ? 1'b0 : n595 ? 1'b0 : 1'b1 : n595 ? 1'b0 : 1'b1 : n1479 ? n705 ? n595 ? 1'b1 : 1'b0 : n595 ? 1'b0 : 1'b1 : n705 ? 1'b1 : n595 ? 1'b0 : 1'b1;
assign n3412 = /* LUT   16 14  2 */ n948 ? n244 ? 1'b0 : n59 ? n525 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n3413 = /* LUT    5 17  0 */ n85 ? n45 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n45 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3414 = /* LUT   14 20  4 */ n865 ? n189 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n189 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n3415 = /* LUT   17 20  3 */ n527 ? 1'b0 : 1'b1;
assign n3416 = /* LUT   19 18  0 */ n35 ? 1'b1 : 1'b0;
assign n3417 = /* LUT   23 15  4 */ n35 ? 1'b1 : 1'b0;
assign n3418 = /* LUT   21 16  2 */ n1579 ? n1663 ? n575 ? 1'b1 : 1'b0 : n1466 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1663 ? 1'b0 : n1466 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n3419 = /* LUT   18 22  4 */ n1025 ? 1'b1 : n1273 ? n641 ? n697 ? 1'b1 : 1'b0 : 1'b1 : n641 ? 1'b0 : 1'b1;
assign n3420 = /* LUT   11 19  0 */ n265 ? 1'b0 : 1'b1;
assign n3421 = /* LUT   22 15  2 */ n238 ? n802 ? n244 ? 1'b0 : n59 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3422 = /* LUT   13 17  6 */ n256 ? 1'b1 : n386 ? 1'b1 : 1'b0;
assign n3423 = /* LUT   18 21  6 */ n731 ? n541 ? n1127 ? n56 ? 1'b1 : 1'b0 : 1'b1 : n1127 ? n56 ? 1'b1 : 1'b0 : 1'b0 : n541 ? 1'b1 : 1'b0;
assign n3424 = /* LUT   19 14  7 */ n1175 ? n1339 ? 1'b1 : n1180 ? 1'b0 : 1'b1 : n1339 ? n1180 ? 1'b1 : 1'b0 : 1'b0;
assign n3425 = /* LUT   16 13  3 */ n770 ? 1'b0 : n42 ? 1'b1 : 1'b0;
assign n3426 = /* LUT    5 18  1 */ n94 ? n53 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n53 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3427 = /* LUT   10 20  7 */ n212 ? 1'b1 : 1'b0;
assign n3428 = /* LUT   13 14  4 */ n42 ? 1'b1 : 1'b0;
assign n3429 = /* LUT   21 15  0 */ n1297 ? n202 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n202 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3430 = /* LUT   20 25  2 */ n44 ? 1'b1 : 1'b0;
assign n3431 = /* LUT   17 21  0 */ n1251 ? 1'b1 : 1'b0;
assign n3432 = /* LUT   19 19  3 */ n35 ? 1'b1 : 1'b0;
assign n3433 = /* LUT   23 12  5 */ n158 ? 1'b1 : 1'b0;
assign n3434 = /* LUT   21 17  1 */ n42 ? 1'b1 : 1'b0;
assign n3435 = /* LUT   18 25  5 */ n725 ? n1281 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1281 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3436 = /* LUT   20 15  2 */ n948 ? n932 ? 1'b0 : n180 ? 1'b0 : n244 ? 1'b0 : 1'b1 : 1'b0;
assign n3437 = /* LUT   11 16  1 */ n357 ? 1'b0 : n489 ? 1'b1 : n342 ? n181 ? 1'b1 : 1'b0 : 1'b1;
assign n3438 = /* LUT   22 14  5 */ n158 ? 1'b1 : 1'b0;
assign n3439 = /* LUT   13 18  7 */ n184 ? 1'b0 : 1'b1;
assign n3440 = /* LUT   15 20  0 */ n836 ? 1'b0 : 1'b1;
assign n3442 = /* LUT   18 20  5 */ n1256 ? n821 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n821 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3443 = /* LUT   23 16  3 */ n42 ? 1'b1 : 1'b0;
assign n3447 = /* LUT   16  7  5 */ n1052 ? n905 ? 1'b0 : 1'b1 : n905 ? 1'b1 : 1'b0;
assign n3448 = /* LUT   19 15  4 */ n1329 ? n1464 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1464 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3449 = /* LUT   16 12  4 */ n591 ? n1071 ? n782 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3450 = /* LUT   10 23  6 */ n218 ? 1'b1 : 1'b0;
assign n3451 = /* LUT   12 12  3 */ io_0_5_1 ? 1'b1 : 1'b0;
assign n3452 = /* LUT   14 22  2 */ n42 ? 1'b1 : 1'b0;
assign n3453 = /* LUT   17 22  1 */ n843 ? 1'b0 : 1'b1;
assign n3454 = /* LUT   19 16  2 */ n44 ? 1'b1 : 1'b0;
assign n3455 = /* LUT   22 10  2 */ n1702 ? n1623 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n1623 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3456 = /* LUT    7 11  1 */ n110 ? n108 ? n109 ? 1'b1 : 1'b0 : n66 ? 1'b1 : 1'b0 : n108 ? n109 ? 1'b1 : 1'b0 : 1'b0;
assign n1673 = /* LUT   21 18  0 */ n575 ? n1180 ? 1'b0 : 1'b1 : n1593 ? n971 ? 1'b0 : n1180 ? 1'b1 : 1'b0 : n971 ? n1180 ? 1'b0 : 1'b1 : 1'b1;
assign n3458 = /* LUT   12 15  7 */ n501 ? 1'b0 : 1'b1;
assign n3459 = /* LUT   18 24  6 */ n218 ? 1'b1 : 1'b0;
assign n3460 = /* LUT   15  7  2 */ n735 ? n906 ? 1'b1 : io_33_1_1 ? 1'b1 : 1'b0 : n906 ? 1'b1 : 1'b0;
assign n1568 = /* LUT   20 14  1 */ n1446 ? n1567 ? n705 ? 1'b0 : 1'b1 : 1'b0 : n1304 ? 1'b1 : n705 ? 1'b1 : 1'b0;
assign n3462 = /* LUT   13 19  0 */ n269 ? 1'b0 : 1'b1;
assign n3463 = /* LUT   18 23  4 */ n49 ? n731 ? n1127 ? 1'b1 : n889 ? 1'b1 : 1'b0 : n889 ? 1'b1 : 1'b0 : n731 ? n1127 ? 1'b0 : n889 ? 1'b1 : 1'b0 : n889 ? 1'b1 : 1'b0;
assign n3464 = /* LUT   14 18  7 */ n834 ? n184 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n184 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n3465 = /* LUT   23 17  4 */ n1729 ? n1746 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1746 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3466 = /* LUT   11 15  3 */ n476 ? n298 ? n32 ? 1'b1 : 1'b0 : n32 ? 1'b0 : 1'b1 : n298 ? n32 ? 1'b0 : 1'b1 : n32 ? 1'b1 : 1'b0;
assign n3467 = /* LUT   14  7  0 */ n739 ? n646 ? 1'b0 : n734 ? 1'b0 : 1'b1 : n646 ? n734 ? 1'b0 : 1'b1 : 1'b0;
assign n3469 = /* LUT   19 12  5 */ n1302 ? n244 ? 1'b0 : n180 ? 1'b0 : n948 ? 1'b1 : 1'b0 : 1'b0;
assign n3470 = /* LUT   16 11  5 */ n158 ? 1'b1 : 1'b0;
assign n3471 = /* LUT   12 19  2 */ n44 ? 1'b1 : 1'b0;
assign n3472 = /* LUT   17 12  7 */ n1161 ? n1152 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1152 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n817  = /* LUT   14 17  3 */ n607 ? n705 ? n816 ? 1'b0 : n595 ? 1'b0 : 1'b1 : n595 ? 1'b0 : 1'b1 : n705 ? n816 ? n595 ? 1'b1 : 1'b0 : 1'b1 : n595 ? 1'b0 : 1'b1;
assign n3474 = /* LUT   17 23  6 */ n989 ? 1'b0 : 1'b1;
assign n3477 = /* LUT   12 14  4 */ n472 ? 1'b0 : 1'b1;
assign n3478 = /* LUT   20 13  0 */ n1295 ? n924 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n924 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3479 = /* LUT   16 23  0 */ io_8_33_1 ? 1'b1 : 1'b0;
assign n3482 = /* LUT   13 20  1 */ n397 ? 1'b0 : 1'b1;
assign n1313 = /* LUT   18 13  2 */ n1293 ? n709 ? n930 ? 1'b0 : 1'b1 : n950 ? 1'b0 : n930 ? 1'b1 : 1'b0 : n709 ? n930 ? 1'b0 : 1'b1 : n950 ? n930 ? 1'b0 : 1'b1 : 1'b1;
assign n3484 = /* LUT   20 19  3 */ n42 ? 1'b1 : 1'b0;
assign n3485 = /* LUT   14 13  6 */ n140 ? 1'b1 : 1'b0;
assign n3486 = /* LUT   23 22  5 */ n218 ? 1'b1 : 1'b0;
assign n1444 = /* LUT   19 13  2 */ n963 ? n1443 ? n575 ? 1'b1 : 1'b0 : n786 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1443 ? 1'b0 : n786 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n3490 = /* LUT   16 10  6 */ n929 ? 1'b1 : 1'b0;
assign n3491 = /* LUT   15 24  1 */ n1027 ? n883 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n883 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3492 = /* LUT   12 18  1 */ n610 ? n485 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n485 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3493 = /* LUT   14 16  0 */ n696 ? n698 ? 1'b0 : n700 ? n699 ? 1'b1 : 1'b0 : 1'b0 : 1'b0;
assign n3494 = /* LUT   17 13  4 */ n1083 ? n1188 ? n709 ? 1'b0 : 1'b1 : n1076 ? 1'b1 : n709 ? 1'b1 : 1'b0 : n1188 ? 1'b0 : n1076 ? 1'b1 : n709 ? 1'b1 : 1'b0;
assign n3495 = /* LUT   21 20  6 */ n140 ? 1'b1 : 1'b0;
assign n3498 = /* LUT    9 17  6 */ n44 ? 1'b1 : 1'b0;
assign n3499 = /* LUT   12 13  5 */ n158 ? 1'b1 : 1'b0;
assign n3500 = /* LUT   18 26  0 */ n1025 ? n28 ? 1'b1 : 1'b0 : n1273 ? n697 ? 1'b1 : n28 ? 1'b1 : 1'b0 : n28 ? 1'b1 : 1'b0;
assign n3501 = /* LUT   16 22  3 */ n731 ? n28 ? 1'b1 : n1127 ? n272 ? 1'b0 : 1'b1 : 1'b0 : n28 ? 1'b1 : 1'b0;
assign n3502 = /* LUT   10 16  4 */ n349 ? n234 ? io_0_25_1 ? 1'b0 : 1'b1 : io_0_25_1 ? 1'b1 : 1'b0 : n234 ? 1'b1 : 1'b0;
assign n3503 = /* LUT   18 12  1 */ n212 ? 1'b1 : 1'b0;
assign n3504 = /* LUT    6 13  3 */ n124 ? 1'b0 : 1'b1;
assign n3505 = /* LUT   20 18  0 */ n1480 ? n1599 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1599 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n774  = /* LUT   14 12  5 */ n157 ? n773 ? 1'b1 : n769 ? io_0_25_1 ? 1'b1 : 1'b0 : 1'b0 : n773 ? 1'b1 : 1'b0;
assign n3507 = /* LUT   11 13  5 */ n218 ? 1'b1 : 1'b0;
assign n3508 = /* LUT   15 25  6 */ n1041 ? n896 ? 1'b0 : n28 ? 1'b0 : 1'b1 : n896 ? n28 ? 1'b0 : 1'b1 : 1'b0;
assign n3509 = /* LUT   12 17  0 */ n356 ? n468 ? 1'b0 ? 1'b1 : 1'b0 : 1'b0 ? 1'b0 : 1'b1 : n468 ? 1'b0 ? 1'b0 : 1'b1 : 1'b0 ? 1'b1 : 1'b0;
assign n3511 = /* LUT   17 14  5 */ n140 ? 1'b1 : 1'b0;
assign n3512 = /* LUT   14 19  1 */ n845 ? n268 ? 1'b0 : n630 ? 1'b0 : 1'b1 : n268 ? n630 ? 1'b0 : 1'b1 : 1'b0;
assign n3513 = /* LUT   17 17  4 */ n212 ? 1'b1 : 1'b0;
assign n3514 = /* LUT   21 21  5 */ n1490 ? n716 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n716 ? n575 ? 1'b1 : 1'b0 : 1'b0;
assign n3515 = /* LUT   16 21  2 */ n35 ? 1'b1 : 1'b0;
assign n3516 = /* LUT   10 19  5 */ n158 ? 1'b1 : 1'b0;
assign n3517 = /* LUT   13 22  3 */ n404 ? 1'b0 : 1'b1;
assign n3518 = /* LUT   18 15  0 */ n780 ? n935 ? n778 ? n943 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n3519 = /* LUT    6 12  0 */ n78 ? 1'b1 : n69 ? n76 ? 1'b1 : n67 ? 1'b0 : 1'b1 : 1'b1;
assign n3520 = /* LUT   20 17  1 */ n159 ? 1'b1 : 1'b0;
assign n3521 = /* LUT   14 15  4 */ n218 ? 1'b1 : 1'b0;
assign n3522 = /* LUT   23 20  7 */ n218 ? 1'b1 : 1'b0;
assign n3523 = /* LUT   19 11  0 */ n159 ? 1'b1 : 1'b0;
assign n3524 = /* LUT   17 15  2 */ n140 ? 1'b1 : 1'b0;
assign n3525 = /* LUT   19 25  1 */ n212 ? 1'b1 : 1'b0;
assign n3528 = /* LUT   22 13  7 */ n1309 ? n1715 ? n575 ? 1'b1 : 1'b0 : n1550 ? 1'b1 : n575 ? 1'b0 : 1'b1 : n1715 ? 1'b0 : n1550 ? 1'b1 : n575 ? 1'b0 : 1'b1;
assign n3529 = /* LUT   11 22  3 */ n140 ? 1'b1 : 1'b0;
assign n3530 = /* LUT   16 15  4 */ n59 ? n1098 ? n244 ? n802 ? 1'b1 : 1'b0 : 1'b0 : 1'b0 : 1'b0;
assign n3531 = /* LUT   16 20  5 */ n540 ? n936 ? n59 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n3532 = /* LUT   15 18  2 */ n44 ? 1'b1 : 1'b0;
assign n3533 = /* LUT   20 16  6 */ n140 ? 1'b1 : 1'b0;
assign n3534 = /* LUT   17 11  7 */ n140 ? 1'b1 : 1'b0;
assign n3535 = /* LUT   11 11  7 */ n422 ? n296 ? 1'b0 : n282 ? 1'b0 : 1'b1 : n296 ? n282 ? 1'b0 : 1'b1 : 1'b0;
assign n3536 = /* LUT   23 14  2 */ n44 ? 1'b1 : 1'b0;
assign n1736 = /* LUT   22 18  0 */ n1670 ? n709 ? n1640 ? 1'b1 : 1'b0 : 1'b0 : n709 ? n1596 ? 1'b1 : 1'b0 : 1'b1;
assign n3538 = /* LUT   21 10  7 */ n1534 ? n1425 ? n1623 ? 1'b0 : n1294 ? 1'b0 : 1'b1 : 1'b0 : 1'b0;
assign n3541 = /* LUT   19 22  0 */ n1510 ? n1389 ? 1'b0 : n1258 ? 1'b0 : 1'b1 : n1389 ? n1258 ? 1'b0 : 1'b1 : 1'b0;
assign n91   = /* CARRY  5 17  5 */ (n49 & 1'b0) | ((n49 | 1'b0) & n90);
assign n1774 = /* CARRY 17 20  6 */ (n1125 & 1'b0) | ((n1125 | 1'b0) & n1828);
assign n1775 = /* CARRY 12 22  5 */ (n515 & n32) | ((n515 | n32) & n1906);
assign n1776 = /* CARRY 11 20  1 */ (n388 & n397) | ((n388 | n397) & n1812);
assign n98   = /* CARRY  5 18  4 */ (n56 & 1'b0) | ((n56 | 1'b0) & n97);
assign n1777 = /* CARRY 17 24  6 */ (n190 & n32) | ((n190 | n32) & n1830);
assign n1778 = /* CARRY 12 21  4 */ (n534 & n183) | ((n534 | n183) & n1814);
assign n458  = /* CARRY 11 14  7 */ (n32 & n438) | ((n32 | n438) & n457);
assign n1779 = /* CARRY 17 22  4 */ (n183 & n1133) | ((n183 | n1133) & n1855);
assign n1708 = /* CARRY 22 10  7 */ (n1540 & 1'b0) | ((n1540 | 1'b0) & n1707);
assign n1780 = /* CARRY 12 15  2 */ (n461 & n325) | ((n461 | n325) & n1832);
assign n1781 = /* CARRY 15 21  4 */ (n873 & n187) | ((n873 | n187) & n1911);
assign n478  = /* CARRY 11 15  4 */ (n32 & n299) | ((n32 | n299) & n477);
assign n511  = /* CARRY 11 18  7 */ (n373 & n184) | ((n373 | n184) & n1816);
assign n1782 = /* CARRY 15 22  6 */ (n190 & n32) | ((n190 | n32) & n1835);
assign n118  = /* CARRY  6 11  5 */ (n72 & 1'b0) | ((n72 | 1'b0) & n117);
assign n1783 = /* CARRY 17 23  3 */ (n1140 & n514) | ((n1140 | n514) & n1913);
assign n1784 = /* CARRY 12 14  1 */ (n443 & n313) | ((n443 | n313) & n1914);
assign n862  = /* CARRY 14 20  0 */ (n398 & 1'b0) | ((n398 | 1'b0) & n852);
assign n287  = /* CARRY 10 10  0 */ (n277 & n194) | ((n277 | n194) & n2014);
assign n1785 = /* CARRY 11 19  4 */ (n379 & n187) | ((n379 | n187) & n1894);
assign n1031 = /* CARRY 15 24  4 */ (n888 & 1'b0) | ((n888 | 1'b0) & n1030);
assign n307  = /* CARRY 10 13  1 */ (n206 & 1'b0) | ((n206 | 1'b0) & n306);
assign n1039 = /* CARRY 15 25  3 */ (n895 & 1'b0) | ((n895 | 1'b0) & n1038);
assign n1786 = /* CARRY 13 18  3 */ (n175 & n130) | ((n175 | n130) & n1819);
assign n1787 = /* CARRY 15 20  4 */ (n857 & n183) | ((n857 | n183) & n1820);
assign n1049 = /* CARRY 16  7  1 */ (n901 & 1'b0) | ((n901 | 1'b0) & n1048);
assign n1788 = /* CARRY 13 19  4 */ (n584 & n617) | ((n584 | n617) & n1873);
assign n831  = /* CARRY 14 18  3 */ (n494 & 1'b0) | ((n494 | 1'b0) & n830);
assign n1789 = /* CARRY 17 18  0 */ (n255 & n979) | ((n255 | n979) & n2063);
assign n335  = /* CARRY 10 15  3 */ (n222 & 1'b0) | ((n222 | 1'b0) & n334);
assign n1790 = /* CARRY 13 23  1 */ (n268 & n32) | ((n268 | n32) & n1917);
assign n416  = /* CARRY 11 11  0 */ (n285 & 1'b0) | ((n285 | 1'b0) & n415);
assign n363  = /* CARRY 10 17  3 */ (n243 & 1'b0) | ((n243 | 1'b0) & n362);
assign n1791 = /* CARRY 13 20  5 */ (n626 & 1'b0) | ((n626 | 1'b0) & n1823);
assign n1792 = /* CARRY 13 24  0 */ (n32 & n398) | ((n32 | n398) & n728);
assign n346  = /* CARRY 10 16  0 */ (n229 & 1'b0) | ((n229 | 1'b0) & n339);
assign n850  = /* CARRY 14 19  5 */ (n515 & 1'b0) | ((n515 | 1'b0) & n849);
assign n1528 = /* CARRY 19 24  2 */ (n1407 & 1'b0) | ((n1407 | 1'b0) & n1527);
assign n1793 = /* CARRY 11 20  4 */ (n391 & n189) | ((n391 | n189) & n1867);
assign n727  = /* CARRY 13 22  7 */ (n639 & n184) | ((n639 | n184) & n1826);
assign n679  = /* CARRY 13 12  1 */ (n560 & 1'b0) | ((n560 | 1'b0) & n678);
assign n1794 = /* CARRY 11 18  2 */ (n368 & n386) | ((n368 | n386) & n1849);
assign n113  = /* CARRY  6 11  0 */ (n67 & 1'b0) | ((n67 | 1'b0) & n112);
assign n87   = /* CARRY  5 17  1 */ (n46 & 1'b0) | ((n46 | 1'b0) & n86);
assign n867  = /* CARRY 14 20  5 */ (n396 & 1'b0) | ((n396 | 1'b0) & n866);
assign n1795 = /* CARRY 17 20  2 */ (n1121 & 1'b0) | ((n1121 | 1'b0) & n1851);
assign n1796 = /* CARRY 11 19  1 */ (n376 & n268) | ((n376 | n268) & n1927);
assign n94   = /* CARRY  5 18  0 */ (n52 & 1'b0) | ((n52 | 1'b0) & n93);
assign n1797 = /* CARRY 13 18  6 */ (n37 & n512) | ((n37 | n512) & n1831);
assign n454  = /* CARRY 11 14  3 */ (n32 & n434) | ((n32 | n434) & n453);
assign n1052 = /* CARRY 16  7  4 */ (n904 & 1'b0) | ((n904 | 1'b0) & n1051);
assign n1798 = /* CARRY 17 22  0 */ (n1129 & n385) | ((n1129 | n385) & n2181);
assign n1704 = /* CARRY 22 10  3 */ (n1624 & 1'b0) | ((n1624 | 1'b0) & n1703);
assign n1799 = /* CARRY 12 15  6 */ (n465 & n329) | ((n465 | n329) & n1856);
assign n1800 = /* CARRY 13 19  1 */ (n186 & n589) | ((n186 | n589) & n1930);
assign n1801 = /* CARRY 15 21  0 */ (n869 & n269) | ((n869 | n269) & n997);
assign n474  = /* CARRY 11 15  0 */ (n32 & n303) | ((n32 | n303) & n458);
assign n1269 = /* CARRY 17 23  7 */ (n513 & n1144) | ((n513 | n1144) & n1931);
assign n1802 = /* CARRY 13 23  6 */ (n32 & n188) | ((n32 | n188) & n1932);
assign n1803 = /* CARRY 12 14  5 */ (n447 & n317) | ((n447 | n317) & n1933);
assign n1804 = /* CARRY 10 10  4 */ (n200 & 1'b0) | ((n200 | 1'b0) & n290);
assign n1805 = /* CARRY 10 17  6 */ (n32 & 1'b0) | ((n32 | 1'b0) & n1861);
assign n1806 = /* CARRY 13 20  0 */ (n621 & 1'b0) | ((n621 | 1'b0) & n717);
assign n1807 = /* CARRY 17 19  4 */ (n877 & n617) | ((n877 | n617) & n1935);
assign n1027 = /* CARRY 15 24  0 */ (n886 & 1'b0) | ((n886 | 1'b0) & n1026);
assign n616  = /* CARRY 12 18  6 */ (n500 & 1'b0) | ((n500 | 1'b0) & n615);
assign n732  = /* CARRY 13 24  7 */ (n526 & n32) | ((n526 | n32) & n1841);
assign n311  = /* CARRY 10 13  5 */ (n209 & 1'b0) | ((n209 | 1'b0) & n310);
assign n351  = /* CARRY 10 16  5 */ (n235 & 1'b0) | ((n235 | 1'b0) & n350);
assign n1043 = /* CARRY 15 25  7 */ (n897 & 1'b0) | ((n897 | 1'b0) & n1042);
assign n604  = /* CARRY 12 17  7 */ (n491 & 1'b0) | ((n491 | 1'b0) & n603);
assign n845  = /* CARRY 14 19  0 */ (n269 & 1'b0) | ((n269 | 1'b0) & n835);
assign n1808 = /* CARRY 13 22  2 */ (n634 & n386) | ((n634 | n386) & n1842);
assign n1809 = /* CARRY 17 18  4 */ (n982 & n605) | ((n982 | n605) & n1843);
assign n339  = /* CARRY 10 15  7 */ (n226 & 1'b0) | ((n226 | 1'b0) & n338);
assign n420  = /* CARRY 11 11  4 */ (n280 & 1'b0) | ((n280 | 1'b0) & n419);
assign n1810 = /* CARRY 12 23  1 */ (n397 & n32) | ((n397 | n32) & n1844);
assign n1514 = /* CARRY 19 22  3 */ (n1392 & 1'b0) | ((n1392 | 1'b0) & n1513);
assign n1811 = /* CARRY 12 22  2 */ (n32 & n516) | ((n32 | n516) & n1920);
assign n1532 = /* CARRY 19 24  6 */ (n796 & 1'b0) | ((n796 | 1'b0) & n1531);
assign n1812 = /* CARRY 11 20  0 */ (n387 & n398) | ((n387 | n398) & n517);
assign n1344 = /* CARRY 18 16  2 */ (n595 & 1'b0) | ((n595 | 1'b0) & n1343);
assign n1813 = /* CARRY 17 24  1 */ (n397 & n32) | ((n397 | n32) & n1846);
assign n1814 = /* CARRY 12 21  3 */ (n494 & n533) | ((n494 | n533) & n1847);
assign n457  = /* CARRY 11 14  6 */ (n32 & n437) | ((n32 | n437) & n456);
assign n1815 = /* CARRY 15 21  5 */ (n874 & n515) | ((n874 | n515) & n1781);
assign n479  = /* CARRY 11 15  5 */ (n32 & n300) | ((n32 | n300) & n478);
assign n1816 = /* CARRY 11 18  6 */ (n372 & n185) | ((n372 | n185) & n1875);
assign n1817 = /* CARRY 15 22  1 */ (n397 & n32) | ((n397 | n32) & n1850);
assign n117  = /* CARRY  6 11  4 */ (n71 & 1'b0) | ((n71 | 1'b0) & n116);
assign n863  = /* CARRY 14 20  1 */ (n397 & 1'b0) | ((n397 | 1'b0) & n862);
assign n288  = /* CARRY 10 10  1 */ (n195 & 1'b0) | ((n195 | 1'b0) & n287);
assign n1818 = /* CARRY 11 19  5 */ (n380 & n515) | ((n380 | n515) & n1785);
assign n306  = /* CARRY 10 13  0 */ (n203 & 1'b0) | ((n203 | 1'b0) & n305);
assign n1819 = /* CARRY 13 18  2 */ (n129 & n142) | ((n129 | n142) & n1853);
assign n1820 = /* CARRY 15 20  3 */ (n856 & n494) | ((n856 | n494) & n1854);
assign n1048 = /* CARRY 16  7  0 */ (n900 & n733) | ((n900 | n733) & n2379);
assign n1821 = /* CARRY 13 19  5 */ (n618 & n585) | ((n618 | n585) & n1788);
assign n832  = /* CARRY 14 18  4 */ (n183 & 1'b0) | ((n183 | 1'b0) & n831);
assign n744  = /* CARRY 14  7  3 */ (n649 & 1'b0) | ((n649 | 1'b0) & n743);
assign n334  = /* CARRY 10 15  2 */ (n221 & 1'b0) | ((n221 | 1'b0) & n333);
assign n1822 = /* CARRY 13 23  2 */ (n32 & n516) | ((n32 | n516) & n1790);
assign n417  = /* CARRY 11 11  1 */ (n283 & 1'b0) | ((n283 | 1'b0) & n416);
assign n362  = /* CARRY 10 17  2 */ (n241 & 1'b0) | ((n241 | 1'b0) & n361);
assign n1823 = /* CARRY 13 20  4 */ (n625 & 1'b0) | ((n625 | 1'b0) & n1839);
assign n1517 = /* CARRY 19 22  6 */ (n1395 & 1'b0) | ((n1395 | 1'b0) & n1516);
assign n1824 = /* CARRY 17 19  0 */ (n267 & n991) | ((n267 | n991) & n1231);
assign n612  = /* CARRY 12 18  2 */ (n486 & 1'b0) | ((n486 | 1'b0) & n611);
assign n1825 = /* CARRY 13 24  3 */ (n527 & n32) | ((n527 | n32) & n1863);
assign n347  = /* CARRY 10 16  1 */ (n231 & 1'b0) | ((n231 | 1'b0) & n346);
assign n600  = /* CARRY 12 17  3 */ (n471 & 1'b0) | ((n471 | 1'b0) & n599);
assign n849  = /* CARRY 14 19  4 */ (n187 & 1'b0) | ((n187 | 1'b0) & n848);
assign n1527 = /* CARRY 19 24  1 */ (n1406 & 1'b0) | ((n1406 | 1'b0) & n1526);
assign n1826 = /* CARRY 13 22  6 */ (n638 & n185) | ((n638 | n185) & n1864);
assign n678  = /* CARRY 13 12  0 */ (n562 & n558) | ((n562 | n558) & n2466);
assign n1827 = /* CARRY 12 23  5 */ (n396 & n32) | ((n396 | n32) & n1865);
assign n92   = /* CARRY  5 17  6 */ (n50 & 1'b0) | ((n50 | 1'b0) & n91);
assign n1828 = /* CARRY 17 20  5 */ (n1124 & 1'b0) | ((n1124 | 1'b0) & n1866);
assign n1829 = /* CARRY 12 22  6 */ (n32 & n188) | ((n32 | n188) & n1775);
assign n101  = /* CARRY  5 18  7 */ (n29 & 1'b0) | ((n29 | 1'b0) & n100);
assign n1830 = /* CARRY 17 24  5 */ (n396 & n32) | ((n396 | n32) & n1868);
assign n631  = /* CARRY 12 21  7 */ (n537 & n184) | ((n537 | n184) & n1869);
assign n1831 = /* CARRY 13 18  5 */ (n177 & n606) | ((n177 | n606) & n1870);
assign n453  = /* CARRY 11 14  2 */ (n32 & n433) | ((n32 | n433) & n452);
assign n102  = /* CARRY  5 19  0 */ (n60 & 1'b0) | ((n60 | 1'b0) & n101);
assign n1263 = /* CARRY 17 22  7 */ (n184 & n1136) | ((n184 | n1136) & n1871);
assign n1705 = /* CARRY 22 10  4 */ (n1294 & 1'b0) | ((n1294 | 1'b0) & n1704);
assign n1832 = /* CARRY 12 15  1 */ (n460 & n324) | ((n460 | n324) & n1872);
assign n1833 = /* CARRY 13 19  2 */ (n582 & n143) | ((n582 | n143) & n1800);
assign n1834 = /* CARRY 15 21  1 */ (n870 & n268) | ((n870 | n268) & n1801);
assign n475  = /* CARRY 11 15  1 */ (n32 & n304) | ((n32 | n304) & n474);
assign n1835 = /* CARRY 15 22  5 */ (n32 & n396) | ((n32 | n396) & n1876);
assign n1836 = /* CARRY 17 23  0 */ (n269 & n1137) | ((n269 | n1137) & n1263);
assign n728  = /* CARRY 13 23  7 */ (n513 & n32) | ((n513 | n32) & n1802);
assign n1837 = /* CARRY 12 14  2 */ (n444 & n314) | ((n444 | n314) & n1784);
assign n1838 = /* CARRY 10 10  5 */ (n32 & 1'b0) | ((n32 | 1'b0) & n1804);
assign n1839 = /* CARRY 13 20  3 */ (n624 & 1'b0) | ((n624 | 1'b0) & n1880);
assign n1840 = /* CARRY 17 19  5 */ (n988 & n618) | ((n988 | n618) & n1807);
assign n1034 = /* CARRY 15 24  7 */ (n891 & 1'b0) | ((n891 | 1'b0) & n1033);
assign n1841 = /* CARRY 13 24  6 */ (n32 & n190) | ((n32 | n190) & n1903);
assign n310  = /* CARRY 10 13  4 */ (n204 & 1'b0) | ((n204 | 1'b0) & n309);
assign n1036 = /* CARRY 15 25  0 */ (n893 & 1'b0) | ((n893 | 1'b0) & n1034);
assign n997  = /* CARRY 15 20  7 */ (n860 & n184) | ((n860 | n184) & n1883);
assign n603  = /* CARRY 12 17  6 */ (n490 & 1'b0) | ((n490 | 1'b0) & n602);
assign n1842 = /* CARRY 13 22  1 */ (n633 & n256) | ((n633 | n256) & n1884);
assign n828  = /* CARRY 14 18  0 */ (n385 & 1'b0) | ((n385 | 1'b0) & n827);
assign n1843 = /* CARRY 17 18  3 */ (n130 & n981) | ((n130 | n981) & n1885);
assign n338  = /* CARRY 10 15  6 */ (n225 & 1'b0) | ((n225 | 1'b0) & n337);
assign n421  = /* CARRY 11 11  5 */ (n281 & 1'b0) | ((n281 | 1'b0) & n420);
assign n1844 = /* CARRY 12 23  0 */ (n32 & n398) | ((n32 | n398) & n640);
assign n1513 = /* CARRY 19 22  2 */ (n1391 & 1'b0) | ((n1391 | 1'b0) & n1512);
assign n1845 = /* CARRY 12 22  3 */ (n514 & n32) | ((n514 | n32) & n1811);
assign n1531 = /* CARRY 19 24  5 */ (n1410 & 1'b0) | ((n1410 | 1'b0) & n1530);
assign n529  = /* CARRY 11 20  7 */ (n394 & n526) | ((n394 | n526) & n1888);
assign n1345 = /* CARRY 18 16  3 */ (n705 & 1'b0) | ((n705 | 1'b0) & n1344);
assign n1846 = /* CARRY 17 24  0 */ (n398 & n32) | ((n398 | n32) & n1269);
assign n1847 = /* CARRY 12 21  2 */ (n386 & n532) | ((n386 | n532) & n1890);
assign n682  = /* CARRY 13 12  4 */ (n568 & 1'b0) | ((n568 | 1'b0) & n681);
assign n1848 = /* CARRY 15 21  6 */ (n875 & n188) | ((n875 | n188) & n1815);
assign n1849 = /* CARRY 11 18  1 */ (n367 & n256) | ((n367 | n256) & n1891);
assign n1850 = /* CARRY 15 22  0 */ (n398 & n32) | ((n398 | n32) & n1006);
assign n116  = /* CARRY  6 11  3 */ (n70 & 1'b0) | ((n70 | 1'b0) & n115);
assign n88   = /* CARRY  5 17  2 */ (n17 & 1'b0) | ((n17 | 1'b0) & n87);
assign n868  = /* CARRY 14 20  6 */ (n190 & 1'b0) | ((n190 | 1'b0) & n867);
assign n1851 = /* CARRY 17 20  1 */ (n1120 & 1'b0) | ((n1120 | 1'b0) & n1893);
assign n289  = /* CARRY 10 10  2 */ (n151 & 1'b0) | ((n151 | 1'b0) & n288);
assign n1852 = /* CARRY 11 19  2 */ (n377 & n516) | ((n377 | n516) & n1796);
assign n97   = /* CARRY  5 18  3 */ (n55 & 1'b0) | ((n55 | 1'b0) & n96);
assign n309  = /* CARRY 10 13  3 */ (n208 & 1'b0) | ((n208 | 1'b0) & n308);
assign n1853 = /* CARRY 13 18  1 */ (n174 & n182) | ((n174 | n182) & n1895);
assign n1854 = /* CARRY 15 20  2 */ (n855 & n386) | ((n855 | n386) & n1896);
assign n1051 = /* CARRY 16  7  3 */ (n903 & 1'b0) | ((n903 | 1'b0) & n1050);
assign n1046 = /* CARRY 15 26  1 */ (n899 & 1'b0) | ((n899 | 1'b0) & n1045);
assign n1855 = /* CARRY 17 22  3 */ (n494 & n1132) | ((n494 | n1132) & n1897);
assign n1701 = /* CARRY 22 10  0 */ (n1425 & n1535) | ((n1425 | n1535) & n2726);
assign n1856 = /* CARRY 12 15  5 */ (n464 & n328) | ((n464 | n328) & n1898);
assign n1857 = /* CARRY 13 19  6 */ (n586 & n524) | ((n586 | n524) & n1821);
assign n833  = /* CARRY 14 18  5 */ (n345 & 1'b0) | ((n345 | 1'b0) & n832);
assign n743  = /* CARRY 14  7  2 */ (n648 & 1'b0) | ((n648 | 1'b0) & n742);
assign n1858 = /* CARRY 17 23  4 */ (n187 & n1141) | ((n187 | n1141) & n1783);
assign n333  = /* CARRY 10 15  1 */ (n220 & 1'b0) | ((n220 | 1'b0) & n332);
assign n1859 = /* CARRY 13 23  3 */ (n514 & n32) | ((n514 | n32) & n1822);
assign n1860 = /* CARRY 12 14  6 */ (n448 & n318) | ((n448 | n318) & n1803);
assign n1861 = /* CARRY 10 17  5 */ (n228 & 1'b0) | ((n228 | 1'b0) & n364);
assign n719  = /* CARRY 13 20  7 */ (n628 & 1'b0) | ((n628 | 1'b0) & n1901);
assign n1862 = /* CARRY 17 19  1 */ (n186 & n992) | ((n186 | n992) & n1824);
assign n1030 = /* CARRY 15 24  3 */ (n887 & 1'b0) | ((n887 | 1'b0) & n1029);
assign n613  = /* CARRY 12 18  3 */ (n487 & 1'b0) | ((n487 | 1'b0) & n612);
assign n1863 = /* CARRY 13 24  2 */ (n32 & n528) | ((n32 | n528) & n1919);
assign n352  = /* CARRY 10 16  6 */ (n236 & 1'b0) | ((n236 | 1'b0) & n351);
assign n1040 = /* CARRY 15 25  4 */ (n541 & 1'b0) | ((n541 | 1'b0) & n1039);
assign n599  = /* CARRY 12 17  2 */ (n470 & 1'b0) | ((n470 | 1'b0) & n598);
assign n848  = /* CARRY 14 19  3 */ (n514 & 1'b0) | ((n514 | 1'b0) & n847);
assign n1526 = /* CARRY 19 24  0 */ (n1405 & 1'b0) | ((n1405 | 1'b0) & n1525);
assign n1864 = /* CARRY 13 22  5 */ (n637 & n345) | ((n637 | n345) & n1904);
assign n1231 = /* CARRY 17 18  7 */ (n983 & n384) | ((n983 | n384) & n1905);
assign n681  = /* CARRY 13 12  3 */ (n567 & 1'b0) | ((n567 | 1'b0) & n680);
assign n1865 = /* CARRY 12 23  4 */ (n32 & n189) | ((n32 | n189) & n1886);
assign n93   = /* CARRY  5 17  7 */ (n27 & 1'b0) | ((n27 | 1'b0) & n92);
assign n1866 = /* CARRY 17 20  4 */ (n1123 & 1'b0) | ((n1123 | 1'b0) & n1926);
assign n640  = /* CARRY 12 22  7 */ (n513 & n32) | ((n513 | n32) & n1829);
assign n1867 = /* CARRY 11 20  3 */ (n390 & n527) | ((n390 | n527) & n1907);
assign n100  = /* CARRY  5 18  6 */ (n58 & 1'b0) | ((n58 | 1'b0) & n99);
assign n1868 = /* CARRY 17 24  4 */ (n189 & n32) | ((n189 | n32) & n1889);
assign n1869 = /* CARRY 12 21  6 */ (n536 & n185) | ((n536 | n185) & n1908);
assign n1870 = /* CARRY 13 18  4 */ (n176 & n605) | ((n176 | n605) & n1786);
assign n456  = /* CARRY 11 14  5 */ (n32 & n436) | ((n32 | n436) & n455);
assign n103  = /* CARRY  5 19  1 */ (n61 & 1'b0) | ((n61 | 1'b0) & n102);
assign n1871 = /* CARRY 17 22  6 */ (n185 & n1135) | ((n185 | n1135) & n1909);
assign n1706 = /* CARRY 22 10  5 */ (n1538 & 1'b0) | ((n1538 | 1'b0) & n1705);
assign n1872 = /* CARRY 12 15  0 */ (n459 & n323) | ((n459 | n323) & n576);
assign n1873 = /* CARRY 13 19  3 */ (n131 & n583) | ((n131 | n583) & n1833);
assign n1874 = /* CARRY 15 21  2 */ (n871 & n516) | ((n871 | n516) & n1834);
assign n480  = /* CARRY 11 15  6 */ (n32 & n301) | ((n32 | n301) & n479);
assign n1875 = /* CARRY 11 18  5 */ (n371 & n345) | ((n371 | n345) & n1912);
assign n1876 = /* CARRY 15 22  4 */ (n189 & n32) | ((n189 | n32) & n1892);
assign n1877 = /* CARRY 17 23  1 */ (n268 & n1138) | ((n268 | n1138) & n1836);
assign n1878 = /* CARRY 12 14  3 */ (n445 & n315) | ((n445 | n315) & n1837);
assign n864  = /* CARRY 14 20  2 */ (n528 & 1'b0) | ((n528 | 1'b0) & n863);
assign n1879 = /* CARRY 10 10  6 */ (n32 & 1'b0) | ((n32 | 1'b0) & n1838);
assign n1880 = /* CARRY 13 20  2 */ (n623 & 1'b0) | ((n623 | 1'b0) & n1934);
assign n1881 = /* CARRY 17 19  6 */ (n989 & n524) | ((n989 | n524) & n1840);
assign n1882 = /* CARRY 11 19  6 */ (n381 & n188) | ((n381 | n188) & n1818);
assign n1033 = /* CARRY 15 24  6 */ (n890 & 1'b0) | ((n890 | 1'b0) & n1032);
assign n614  = /* CARRY 12 18  4 */ (n499 & 1'b0) | ((n499 | 1'b0) & n613);
assign n1037 = /* CARRY 15 25  1 */ (n892 & 1'b0) | ((n892 | 1'b0) & n1036);
assign n1883 = /* CARRY 15 20  6 */ (n185 & n859) | ((n185 | n859) & n1915);
assign n602  = /* CARRY 12 17  5 */ (n473 & 1'b0) | ((n473 | 1'b0) & n601);
assign n1884 = /* CARRY 13 22  0 */ (n385 & n632) | ((n385 | n632) & n2939);
assign n829  = /* CARRY 14 18  1 */ (n256 & 1'b0) | ((n256 | 1'b0) & n828);
assign n1885 = /* CARRY 17 18  2 */ (n142 & n980) | ((n142 | n980) & n1916);
assign n337  = /* CARRY 10 15  5 */ (n224 & 1'b0) | ((n224 | 1'b0) & n336);
assign n418  = /* CARRY 11 11  2 */ (n294 & 1'b0) | ((n294 | 1'b0) & n417);
assign n361  = /* CARRY 10 17  1 */ (n240 & 1'b0) | ((n240 | 1'b0) & n360);
assign n1886 = /* CARRY 12 23  3 */ (n527 & n32) | ((n527 | n32) & n1918);
assign n1516 = /* CARRY 19 22  5 */ (n1394 & 1'b0) | ((n1394 | 1'b0) & n1515);
assign n348  = /* CARRY 10 16  2 */ (n232 & 1'b0) | ((n232 | 1'b0) & n347);
assign n1887 = /* CARRY 12 22  0 */ (n32 & n269) | ((n32 | n269) & n631);
assign n852  = /* CARRY 14 19  7 */ (n513 & 1'b0) | ((n513 | 1'b0) & n851);
assign n1530 = /* CARRY 19 24  4 */ (n1409 & 1'b0) | ((n1409 | 1'b0) & n1529);
assign n1888 = /* CARRY 11 20  6 */ (n393 & n190) | ((n393 | n190) & n1921);
assign n1342 = /* CARRY 18 16  0 */ (n575 & n930) | ((n575 | n930) & n3003);
assign n1889 = /* CARRY 17 24  3 */ (n32 & n527) | ((n32 | n527) & n1922);
assign n1890 = /* CARRY 12 21  1 */ (n531 & n256) | ((n531 | n256) & n1923);
assign n1006 = /* CARRY 15 21  7 */ (n876 & n513) | ((n876 | n513) & n1848);
assign n1891 = /* CARRY 11 18  0 */ (n366 & n385) | ((n366 | n385) & n3034);
assign n1892 = /* CARRY 15 22  3 */ (n527 & n32) | ((n527 | n32) & n1925);
assign n115  = /* CARRY  6 11  2 */ (n69 & 1'b0) | ((n69 | 1'b0) & n114);
assign n89   = /* CARRY  5 17  3 */ (n47 & 1'b0) | ((n47 | 1'b0) & n88);
assign n1893 = /* CARRY 17 20  0 */ (n1119 & 1'b0) | ((n1119 | 1'b0) & n1244);
assign n290  = /* CARRY 10 10  3 */ (n152 & 1'b0) | ((n152 | 1'b0) & n289);
assign n1894 = /* CARRY 11 19  3 */ (n378 & n514) | ((n378 | n514) & n1852);
assign n96   = /* CARRY  5 18  2 */ (n54 & 1'b0) | ((n54 | 1'b0) & n95);
assign n308  = /* CARRY 10 13  2 */ (n207 & 1'b0) | ((n207 | 1'b0) & n307);
assign n1895 = /* CARRY 13 18  0 */ (n173 & n255) | ((n173 | n255) & n3082);
assign n1896 = /* CARRY 15 20  1 */ (n854 & n256) | ((n854 | n256) & n1928);
assign n452  = /* CARRY 11 14  1 */ (n32 & n432) | ((n32 | n432) & n451);
assign n1050 = /* CARRY 16  7  2 */ (n902 & 1'b0) | ((n902 | 1'b0) & n1049);
assign n1045 = /* CARRY 15 26  0 */ (n898 & 1'b0) | ((n898 | 1'b0) & n1043);
assign n1897 = /* CARRY 17 22  2 */ (n386 & n1131) | ((n386 | n1131) & n1929);
assign n1702 = /* CARRY 22 10  1 */ (n1622 & 1'b0) | ((n1622 | 1'b0) & n1701);
assign n1898 = /* CARRY 12 15  4 */ (n463 & n327) | ((n463 | n327) & n1910);
assign n717  = /* CARRY 13 19  7 */ (n395 & n587) | ((n395 | n587) & n1857);
assign n834  = /* CARRY 14 18  6 */ (n185 & 1'b0) | ((n185 | 1'b0) & n833);
assign n476  = /* CARRY 11 15  2 */ (n32 & n297) | ((n32 | n297) & n475);
assign n742  = /* CARRY 14  7  1 */ (n647 & 1'b0) | ((n647 | 1'b0) & n741);
assign n1899 = /* CARRY 17 23  5 */ (n515 & n1142) | ((n515 | n1142) & n1858);
assign n332  = /* CARRY 10 15  0 */ (n213 & n214) | ((n213 | n214) & n3111);
assign n1900 = /* CARRY 13 23  4 */ (n32 & n187) | ((n32 | n187) & n1859);
assign n576  = /* CARRY 12 14  7 */ (n449 & n319) | ((n449 | n319) & n1860);
assign n364  = /* CARRY 10 17  4 */ (n227 & 1'b0) | ((n227 | 1'b0) & n363);
assign n1901 = /* CARRY 13 20  6 */ (n627 & 1'b0) | ((n627 | 1'b0) & n1791);
assign n1902 = /* CARRY 17 19  2 */ (n143 & n878) | ((n143 | n878) & n1862);
assign n1029 = /* CARRY 15 24  2 */ (n884 & 1'b0) | ((n884 | 1'b0) & n1028);
assign n610  = /* CARRY 12 18  0 */ (n484 & 1'b0) | ((n484 | 1'b0) & n604);
assign n1903 = /* CARRY 13 24  5 */ (n396 & n32) | ((n396 | n32) & n1936);
assign n353  = /* CARRY 10 16  7 */ (n237 & 1'b0) | ((n237 | 1'b0) & n352);
assign n1041 = /* CARRY 15 25  5 */ (n885 & 1'b0) | ((n885 | 1'b0) & n1040);
assign n598  = /* CARRY 12 17  1 */ (n469 & 1'b0) | ((n469 | 1'b0) & n597);
assign n847  = /* CARRY 14 19  2 */ (n516 & 1'b0) | ((n516 | 1'b0) & n846);
assign n1904 = /* CARRY 13 22  4 */ (n183 & n636) | ((n183 | n636) & n1937);
assign n1905 = /* CARRY 17 18  6 */ (n861 & n512) | ((n861 | n512) & n1938);
assign n680  = /* CARRY 13 12  2 */ (n559 & 1'b0) | ((n559 | 1'b0) & n679);
assign n422  = /* CARRY 11 11  6 */ (n295 & 1'b0) | ((n295 | 1'b0) & n421);
assign n642  = /* CARRY 12 23  7 */ (n526 & n32) | ((n526 | n32) & n1939);
assign n1512 = /* CARRY 19 22  1 */ (n1390 & 1'b0) | ((n1390 | 1'b0) & n1511);
assign n90   = /* CARRY  5 17  4 */ (n48 & 1'b0) | ((n48 | 1'b0) & n89);
assign n1251 = /* CARRY 17 20  7 */ (n1126 & 1'b0) | ((n1126 | 1'b0) & n1774);
assign n1906 = /* CARRY 12 22  4 */ (n32 & n187) | ((n32 | n187) & n1845);
assign n1907 = /* CARRY 11 20  2 */ (n389 & n528) | ((n389 | n528) & n1776);
assign n99   = /* CARRY  5 18  5 */ (n57 & 1'b0) | ((n57 | 1'b0) & n98);
assign n1274 = /* CARRY 17 24  7 */ (n526 & n32) | ((n526 | n32) & n1777);
assign n1908 = /* CARRY 12 21  5 */ (n535 & n345) | ((n535 | n345) & n1778);
assign n455  = /* CARRY 11 14  4 */ (n32 & n435) | ((n32 | n435) & n454);
assign n1909 = /* CARRY 17 22  5 */ (n345 & n1134) | ((n345 | n1134) & n1779);
assign n1707 = /* CARRY 22 10  6 */ (n1626 & 1'b0) | ((n1626 | 1'b0) & n1706);
assign n1910 = /* CARRY 12 15  3 */ (n462 & n326) | ((n462 | n326) & n1780);
assign n1911 = /* CARRY 15 21  3 */ (n872 & n514) | ((n872 | n514) & n1874);
assign n745  = /* CARRY 14  7  4 */ (n650 & 1'b0) | ((n650 | 1'b0) & n744);
assign n1912 = /* CARRY 11 18  4 */ (n370 & n183) | ((n370 | n183) & n1924);
assign n1013 = /* CARRY 15 22  7 */ (n32 & n526) | ((n32 | n526) & n1782);
assign n119  = /* CARRY  6 11  6 */ (n73 & 1'b0) | ((n73 | 1'b0) & n118);
assign n1913 = /* CARRY 17 23  2 */ (n516 & n1139) | ((n516 | n1139) & n1877);
assign n1914 = /* CARRY 12 14  0 */ (n442 & n572) | ((n442 | n572) & n3267);
assign n865  = /* CARRY 14 20  3 */ (n527 & 1'b0) | ((n527 | 1'b0) & n864);
assign n291  = /* CARRY 10 10  7 */ (n32 & 1'b0) | ((n32 | 1'b0) & n1879);
assign n1244 = /* CARRY 17 19  7 */ (n990 & n395) | ((n990 | n395) & n1881);
assign n517  = /* CARRY 11 19  7 */ (n382 & n513) | ((n382 | n513) & n1882);
assign n1032 = /* CARRY 15 24  5 */ (n889 & 1'b0) | ((n889 | 1'b0) & n1031);
assign n615  = /* CARRY 12 18  5 */ (n488 & 1'b0) | ((n488 | 1'b0) & n614);
assign n312  = /* CARRY 10 13  6 */ (n210 & 1'b0) | ((n210 | 1'b0) & n311);
assign n1038 = /* CARRY 15 25  2 */ (n894 & 1'b0) | ((n894 | 1'b0) & n1037);
assign n1915 = /* CARRY 15 20  5 */ (n858 & n345) | ((n858 | n345) & n1787);
assign n601  = /* CARRY 12 17  4 */ (n472 & 1'b0) | ((n472 | 1'b0) & n600);
assign n830  = /* CARRY 14 18  2 */ (n386 & 1'b0) | ((n386 | 1'b0) & n829);
assign n1916 = /* CARRY 17 18  1 */ (n182 & n843) | ((n182 | n843) & n1789);
assign n336  = /* CARRY 10 15  4 */ (n223 & 1'b0) | ((n223 | 1'b0) & n335);
assign n1917 = /* CARRY 13 23  0 */ (n32 & n269) | ((n32 | n269) & n727);
assign n419  = /* CARRY 11 11  3 */ (n286 & 1'b0) | ((n286 | 1'b0) & n418);
assign n360  = /* CARRY 10 17  0 */ (n242 & 1'b0) | ((n242 | 1'b0) & n353);
assign n1918 = /* CARRY 12 23  2 */ (n32 & n528) | ((n32 | n528) & n1810);
assign n1515 = /* CARRY 19 22  4 */ (n1393 & 1'b0) | ((n1393 | 1'b0) & n1514);
assign n1919 = /* CARRY 13 24  1 */ (n397 & n32) | ((n397 | n32) & n1792);
assign n349  = /* CARRY 10 16  3 */ (n233 & 1'b0) | ((n233 | 1'b0) & n348);
assign n1920 = /* CARRY 12 22  1 */ (n268 & n32) | ((n268 | n32) & n1887);
assign n851  = /* CARRY 14 19  6 */ (n188 & 1'b0) | ((n188 | 1'b0) & n850);
assign n1529 = /* CARRY 19 24  3 */ (n1408 & 1'b0) | ((n1408 | 1'b0) & n1528);
assign n1921 = /* CARRY 11 20  5 */ (n392 & n396) | ((n392 | n396) & n1793);
assign n1343 = /* CARRY 18 16  1 */ (n709 & 1'b0) | ((n709 | 1'b0) & n1342);
assign n1922 = /* CARRY 17 24  2 */ (n528 & n32) | ((n528 | n32) & n1813);
assign n1923 = /* CARRY 12 21  0 */ (n530 & n385) | ((n530 | n385) & n3378);
assign n1924 = /* CARRY 11 18  3 */ (n369 & n494) | ((n369 | n494) & n1794);
assign n1925 = /* CARRY 15 22  2 */ (n528 & n32) | ((n528 | n32) & n1817);
assign n114  = /* CARRY  6 11  1 */ (n68 & 1'b0) | ((n68 | 1'b0) & n113);
assign n86   = /* CARRY  5 17  0 */ (n45 & 1'b0) | ((n45 | 1'b0) & n85);
assign n866  = /* CARRY 14 20  4 */ (n189 & 1'b0) | ((n189 | 1'b0) & n865);
assign n1926 = /* CARRY 17 20  3 */ (n1122 & 1'b0) | ((n1122 | 1'b0) & n1795);
assign n1927 = /* CARRY 11 19  0 */ (n375 & n269) | ((n375 | n269) & n511);
assign n95   = /* CARRY  5 18  1 */ (n53 & 1'b0) | ((n53 | 1'b0) & n94);
assign n715  = /* CARRY 13 18  7 */ (n178 & n384) | ((n178 | n384) & n1797);
assign n1928 = /* CARRY 15 20  0 */ (n853 & n385) | ((n853 | n385) & n3441);
assign n451  = /* CARRY 11 14  0 */ (1'b0 & n431) | ((1'b0 | n431) & n3446);
assign n1929 = /* CARRY 17 22  1 */ (n1130 & n256) | ((n1130 | n256) & n1798);
assign n1703 = /* CARRY 22 10  2 */ (n1623 & 1'b0) | ((n1623 | 1'b0) & n1702);
assign n581  = /* CARRY 12 15  7 */ (n466 & n330) | ((n466 | n330) & n1799);
assign n1930 = /* CARRY 13 19  0 */ (n588 & n267) | ((n588 | n267) & n715);
assign n835  = /* CARRY 14 18  7 */ (n184 & 1'b0) | ((n184 | 1'b0) & n834);
assign n477  = /* CARRY 11 15  3 */ (n32 & n298) | ((n32 | n298) & n476);
assign n741  = /* CARRY 14  7  0 */ (n646 & n739) | ((n646 | n739) & n3468);
assign n1931 = /* CARRY 17 23  6 */ (n188 & n1143) | ((n188 | n1143) & n1899);
assign n1932 = /* CARRY 13 23  5 */ (n515 & n32) | ((n515 | n32) & n1900);
assign n1933 = /* CARRY 12 14  4 */ (n446 & n316) | ((n446 | n316) & n1878);
assign n365  = /* CARRY 10 17  7 */ (1'b0 & n32) | ((1'b0 | n32) & n1805);
assign n1934 = /* CARRY 13 20  1 */ (n622 & 1'b0) | ((n622 | 1'b0) & n1806);
assign n1935 = /* CARRY 17 19  3 */ (n131 & n987) | ((n131 | n987) & n1902);
assign n1028 = /* CARRY 15 24  1 */ (n883 & 1'b0) | ((n883 | 1'b0) & n1027);
assign n611  = /* CARRY 12 18  1 */ (n485 & 1'b0) | ((n485 | 1'b0) & n610);
assign n1936 = /* CARRY 13 24  4 */ (n32 & n189) | ((n32 | n189) & n1825);
assign n350  = /* CARRY 10 16  4 */ (n234 & 1'b0) | ((n234 | 1'b0) & n349);
assign n1042 = /* CARRY 15 25  6 */ (n896 & 1'b0) | ((n896 | 1'b0) & n1041);
assign n597  = /* CARRY 12 17  0 */ (n468 & n356) | ((n468 | n356) & n3510);
assign n846  = /* CARRY 14 19  1 */ (n268 & 1'b0) | ((n268 | 1'b0) & n845);
assign n1937 = /* CARRY 13 22  3 */ (n635 & n494) | ((n635 | n494) & n1808);
assign n1938 = /* CARRY 17 18  5 */ (n844 & n606) | ((n844 | n606) & n1809);
assign n1939 = /* CARRY 12 23  6 */ (n32 & n190) | ((n32 | n190) & n1827);
assign n1511 = /* CARRY 19 22  0 */ (n1389 & 1'b0) | ((n1389 | 1'b0) & n1510);
/* FF 16 16  2 */ always @(posedge n3, posedge n5) if (n5) n962 <= 1'b0; else if (n799) n962 <= n1940;
/* FF 22 12  4 */ always @(posedge n3, posedge n5) if (n5) n1636 <= 1'b0; else if (n1077) n1636 <= n1941;
/* FF 15 13  0 */ assign n1942 = n945;
/* FF 20 20  3 */ always @(posedge n3, posedge n5) if (n5) n721 <= 1'b0; else if (n996) n721 <= n1943;
/* FF 16 14  7 */ assign n949 = n1944;
/* FF  5 17  5 */ always @(posedge n3, posedge n5) if (n5) n49 <= 1'b0; else if (n4) n49 <= n1945;
/* FF 16 19  4 */ always @(posedge n3, posedge n5) if (n5) n989 <= 1'b0; else if (n801) n989 <= n1946;
/* FF 15 19  1 */ always @(posedge n3, posedge n5) if (n5) n837 <= 1'b0; else if (n629) n837 <= n1947;
/* FF 17 20  6 */ assign n1125 = n1948;
/* FF 23 15  1 */ always @(posedge n3, posedge n5) if (n5) n1340 <= 1'b0; else if (n1654) n1340 <= n1949;
/* FF 24 16  1 */ always @(posedge n3, posedge n5) if (n5) n1743 <= 1'b0; else if (n619) n1743 <= n1950;
/* FF  7 16  7 */ always @(posedge n3, posedge n5) if (n5) n51 <= 1'b0; else if (1'b1) n51 <= n1951;
/* FF 21 11  0 */ always @(posedge n3, posedge n5) if (n5) n1177 <= 1'b0; else if (n1631) n1177 <= n1952;
/* FF 12 22  5 */ assign n1953 = n1954;
/* FF 19 23  3 */ always @(posedge n3, posedge n5) if (n5) n1401 <= 1'b0; else if (1'b1) n1401 <= n1955;
/* FF 10  9  5 */ always @(posedge n1, posedge n5) if (n5) n152 <= 1'b0; else if (1'b1) n152 <= n1956;
/* FF 22 15  5 */ assign n1654 = n1957;
/* FF 20 11  2 */ always @(posedge n3, posedge n5) if (n5) n1429 <= 1'b0; else if (n1199) n1429 <= n1958;
/* FF 19 24  7 */ always @(posedge n3, posedge n5) if (n5) n797 <= 1'b0; else if (n1025) n797 <= n1959;
/* FF 11 20  1 */ assign n388 = n1960;
/* FF 16 13  6 */ assign n937 = n1079;
/* FF  5 18  4 */ always @(posedge n3, posedge n5) if (n5) n56 <= 1'b0; else if (n4) n56 <= n1961;
/* FF 16 18  7 */ always @(posedge n3, posedge n5) if (n5) n983 <= 1'b1; else if (n800) n983 <= n1962;
/* FF 10 20  0 */ always @(posedge n3, posedge n5) if (n5) n259 <= 1'b1; else if (n144) n259 <= n1963;
/* FF 21 15  5 */ always @(posedge n3, posedge n5) if (n5) n1574 <= 1'b0; else if (n933) n1574 <= n1964;
/* FF 20 22  4 */ assign n641 = n1965;
/* FF 17 21  5 */ assign n1128 = n1966;
/* FF 17 24  6 */ assign n1967 = n1968;
/* FF 23 12  0 */ always @(posedge n3) if (n1301) n960 <= 1'b0 ? 1'b0 : n1969;
/* FF 24 15  0 */ always @(posedge n3, posedge n5) if (n5) n171 <= 1'b0; else if (n958) n171 <= n1970;
/* FF 21 12  1 */ always @(posedge n3, posedge n5) if (n5) n1546 <= 1'b0; else if (n1186) n1546 <= n1971;
/* FF 12 21  4 */ assign n534 = n1972;
/* FF 17 10  1 */ always @(posedge n1, posedge n5) if (n5) n564 <= 1'b0; else if (n8) n564 <= n1973;
/* FF 19 20  2 */ always @(posedge n3, posedge n5) if (n5) n1378 <= 1'b0; else if (1'b1) n1378 <= n1974;
/* FF 22 14  2 */ always @(posedge n3, posedge n5) if (n5) n1646 <= 1'b0; else if (n1651) n1646 <= n1975;
/* FF 23 16  6 */ always @(posedge n3, posedge n5) if (n5) n1485 <= 1'b0; else if (n1653) n1485 <= n1976;
/* FF 11 14  7 */ assign n319 = n1977;
/* FF 16 12  1 */ always @(posedge n3, posedge n5) if (n5) n440 <= 1'b0; else if (n321) n440 <= n1978;
/* FF 16 17  6 */ always @(posedge n3, posedge n5) if (n5) n970 <= 1'b0; else if (n702) n970 <= n1979;
/* FF 13 15  0 */ always @(posedge n3) if (io_0_25_1) n577 <= 1'b0 ? 1'b0 : n1980;
/* FF 15 17  7 */ always @(posedge n3, posedge n5) if (n5) n813 <= 1'b0; else if (n609) n813 <= n1981;
/* FF 20 24  2 */ assign n1523 = n1982;
/* FF 20 21  5 */ always @(posedge n3, posedge n5) if (n5) n1498 <= 1'b0; else if (n1012) n1498 <= n1983;
/* FF 17 22  4 */ assign n1133 = n1984;
/* FF 24 14  3 */ always @(posedge n3, posedge n5) if (n5) n1583 <= 1'b0; else if (n467) n1583 <= n1985;
/* FF 22 10  7 */ always @(posedge n1, posedge n5) if (n5) n1540 <= 1'b0; else if (1'b1) n1540 <= n1986;
/* FF 21 13  2 */ assign n1987 = n1644;
/* FF 12 15  2 */ assign n461 = n1988;
/* FF 19 21  5 */ always @(posedge n3, posedge n5) if (n5) n1283 <= 1'b1; else if (n1145) n1283 <= n1989;
/* FF 11 17  3 */ assign n354 = n496;
/* FF 16  8  6 */ always @(posedge n1, posedge n5) if (n5) n909 <= 1'b0; else if (n8) n909 <= n1990;
/* FF 24 17  7 */ always @(posedge n3, posedge n5) if (n5) n644 <= 1'b0; else if (n1454) n644 <= n1991;
/* FF 15 21  4 */ assign n873 = n1992;
/* FF 23 17  1 */ assign n1993 = n1745;
/* FF 11 15  4 */ assign n327 = n1994;
/* FF 11 18  7 */ assign n373 = n1995;
/* FF 16 11  0 */ always @(posedge n3, posedge n5) if (n5) n923 <= 1'b0; else if (n938) n923 <= n1996;
/* FF 13 16  1 */ always @(posedge n3, posedge n5) if (n5) n583 <= 1'b0; else if (n492) n583 <= n1997;
/* FF 15 22  6 */ assign n1998 = n1999;
/* FF 18  9  2 */ always @(posedge n3, posedge n5) if (n5) n915 <= 1'b0; else if (n215) n915 <= n2000;
/* FF  6 11  5 */ always @(posedge n1, posedge n5) if (n5) n72 <= 1'b0; else if (1'b1) n72 <= n2001;
/* FF 12 24  0 */ assign n542 = n2002;
/* FF 17 23  3 */ assign n1140 = n2003;
/* FF 19 17  2 */ always @(posedge n1, posedge n5) if (n5) n929 <= 1'b0; else if (n8) n929 <= n2004;
/* FF 22 21  5 */ always @(posedge n3, posedge n5) if (n5) n1362 <= 1'b0; else if (n1652) n1362 <= n2005;
/* FF 24 13  2 */ always @(posedge n3, posedge n5) if (n5) n1111 <= 1'b0; else if (n805) n1111 <= n2006;
/* FF 21 14  3 */ assign n2007 = n1649;
/* FF  9 16  0 */ assign n166 = n2008;
/* FF 12 14  1 */ assign n443 = n2009;
/* FF 14 20  0 */ always @(posedge n3, posedge n5) if (n5) n398 <= 1'b0; else if (1'b1) n398 <= n2010;
/* FF 19 18  4 */ assign n2011 = n1489;
/* FF 10 10  0 */ assign n2012 = n2013;
/* FF 16 23  7 */ always @(posedge n3, posedge n5) if (n5) n104 <= 1'b0; else if (n1010) n104 <= n2015;
/* FF 15 10  5 */ always @(posedge n1, posedge n5) if (n5) n672 <= 1'b1; else if (1'b1) n672 <= n2016;
/* FF 20 19  6 */ always @(posedge n3, posedge n5) if (n5) n1373 <= 1'b0; else if (n803) n1373 <= n2017;
/* FF 18 22  0 */ assign n881 = n2018;
/* FF 11 12  5 */ always @(posedge n3, posedge n5) if (n5) n158 <= 1'b0; else if (n26) n158 <= n2019;
/* FF 11 19  4 */ assign n379 = n2020;
/* FF 16 10  3 */ always @(posedge n1, posedge n5) if (n5) n920 <= 1'b0; else if (n672) n920 <= n2021;
/* FF  9 12  2 */ assign n2022 = n205;
/* FF 15 24  4 */ always @(posedge n3, posedge n5) if (n5) n888 <= 1'b0; else if (n2) n888 <= n2023;
/* FF 13 17  2 */ assign n2024 = n710;
/* FF 17 16  2 */ assign n2025 = n1212;
/* FF 19 14  3 */ assign n2026 = n1451;
/* FF 22 20  6 */ assign n1687 = n2027;
/* FF 16 24  3 */ always @(posedge n3, posedge n5) if (n5) n274 <= 1'b0; else if (n1010) n274 <= n2028;
/* FF 12 13  0 */ always @(posedge n3, posedge n5) if (n5) n431 <= 1'b0; else if (n573) n431 <= n2029;
/* FF 20 12  4 */ always @(posedge n3, posedge n5) if (n5) n1308 <= 1'b0; else if (n1299) n1308 <= n2030;
/* FF 10 13  1 */ always @(posedge n1, posedge n5) if (n5) n206 <= 1'b0; else if (n138) n206 <= n2031;
/* FF 16 22  4 */ assign n1010 = n2032;
/* FF 15 11  6 */ always @(posedge n1, posedge n5) if (n5) n765 <= 1'b0; else if (1'b1) n765 <= n2033;
/* FF 20 18  5 */ assign n1481 = n2034;
/* FF 20 15  6 */ assign n805 = n2035;
/* FF 11 13  2 */ always @(posedge n3, posedge n5) if (n5) n299 <= 1'b0; else if (n441) n299 <= n2036;
/* FF 11 16  5 */ assign n342 = n2037;
/* FF  9 13  1 */ always @(posedge n3, posedge n5) if (n5) n44 <= 1'b0; else if (n26) n44 <= n2038;
/* FF 15 25  3 */ always @(posedge n3, posedge n5) if (n5) n895 <= 1'b0; else if (n2) n895 <= n2039;
/* FF 13 18  3 */ assign n130 = n2040;
/* FF 18 11  0 */ always @(posedge n3, posedge n5) if (n5) n1159 <= 1'b0; else if (n1179) n1159 <= n2041;
/* FF 15 20  4 */ assign n857 = n2042;
/* FF 17 17  1 */ assign n2043 = n1220;
/* FF 16  7  1 */ always @(negedge io_0_6_1, posedge n5) if (n5) n901 <= 1'b0; else if (1'b1) n901 <= n2044;
/* FF 19 15  0 */ always @(posedge n3, posedge n5) if (n5) n1327 <= 1'b0; else if (n619) n1327 <= n2045;
/* FF 22 23  7 */ always @(posedge n3, posedge n5) if (n5) n1419 <= 1'b0; else if (n1656) n1419 <= n2046;
/* FF  9 18  2 */ always @(posedge n3, posedge n5) if (n5) n37 <= 1'b1; else if (n172) n37 <= n2047;
/* FF 11  9  7 */ always @(posedge n1, posedge n5) if (n5) n151 <= 1'b0; else if (1'b1) n151 <= n2048;
/* FF 19 16  6 */ always @(posedge n3, posedge n5) if (n5) n1339 <= 1'b0; else if (n949) n1339 <= n2049;
/* FF 16 21  5 */ always @(posedge n3, posedge n5) if (n5) n1003 <= 1'b0; else if (n995) n1003 <= n2050;
/* FF 15  8  7 */ assign n645 = n2051;
/* FF  6 12  5 */ always @(posedge n1, posedge n5) if (n5) n79 <= 1'b0; else if (1'b1) n79 <= n2052;
/* FF 15  7  6 */ assign n739 = n2053;
/* FF 18 24  2 */ assign n1271 = n2054;
/* FF 20 17  4 */ assign n1471 = n2055;
/* FF 20 14  5 */ assign n1446 = n2056;
/* FF 23 20  2 */ always @(posedge n3, posedge n5) if (n5) n1699 <= 1'b0; else if (n1655) n1699 <= n2057;
/* FF 11 10  3 */ assign n284 = n2058;
/* FF 13 19  4 */ assign n617 = n2059;
/* FF 14 18  3 */ always @(posedge n3, posedge n5) if (n5) n494 <= 1'b0; else if (1'b1) n494 <= n2060;
/* FF 17 18  0 */ assign n2061 = n2062;
/* FF 19 12  1 */ assign n1298 = n2064;
/* FF 17 12  3 */ assign n1065 = n2065;
/* FF 10 15  3 */ always @(posedge n1) if (1'b1) n222 <= n7 ? 1'b0 : n2066;
/* FF 16 20  2 */ assign n826 = n2067;
/* FF 13 23  1 */ assign n2068 = n2069;
/* FF 15  9  0 */ always @(posedge n3, posedge n5) if (n5) n652 <= 1'b0; else if (1'b1) n652 <= n2070;
/* FF 18 14  4 */ assign n2071 = n1326;
/* FF 20 16  3 */ always @(posedge n3, posedge n5) if (n5) n1467 <= 1'b0; else if (n1455) n1467 <= n2072;
/* FF 20 13  4 */ assign n1438 = n2073;
/* FF 11 11  0 */ assign n292 = n2074;
/* FF 22 18  5 */ assign n2075 = n1739;
/* FF 10 17  3 */ always @(posedge n1) if (1'b1) n243 <= n7 ? 1'b0 : n2076;
/* FF  9 15  7 */ assign n164 = n2077;
/* FF 13 20  5 */ assign n626 = n2078;
/* FF 18 13  6 */ assign n2079 = n1315;
/* FF 14 13  2 */ always @(posedge n3, posedge n5) if (n5) n684 <= 1'b0; else if (n690) n684 <= n2080;
/* FF 19 22  7 */ always @(posedge n3, posedge n5) if (n5) n1396 <= 1'b0; else if (1'b1) n1396 <= n2081;
/* FF 19 13  6 */ assign n1306 = n2082;
/* FF 23 11  1 */ always @(posedge n3, posedge n5) if (n5) n1556 <= 1'b0; else if (n938) n1556 <= n2083;
/* FF 22 17  1 */ always @(posedge n1, posedge n5) if (n5) n1056 <= 1'b0; else if (n8) n1056 <= n2084;
/* FF 16 16  7 */ always @(posedge n3, posedge n5) if (n5) n968 <= 1'b0; else if (n799) n968 <= n2085;
/* FF 15 13  5 */ assign n777 = n2086;
/* FF 17 13  0 */ always @(posedge n3, posedge n5) if (n5) n1073 <= 1'b0; else if (n596) n1073 <= n2087;
/* FF 14 16  4 */ assign n2088 = n807;
/* FF 16 19  3 */ always @(posedge n3, posedge n5) if (n5) n988 <= 1'b1; else if (n801) n988 <= n2089;
/* FF 13 24  0 */ assign n2090 = n2091;
/* FF 15 14  1 */ assign n781 = n956;
/* FF 18 17  5 */ assign n2092 = n1354;
/* FF 20 23  2 */ always @(posedge n3) if (n688) n1518 <= 1'b0 ? 1'b0 : n2093;
/* FF 10 16  0 */ always @(posedge n1) if (1'b1) n229 <= n7 ? 1'b0 : n2094;
/* FF 13 10  7 */ always @(posedge n1, posedge n5) if (n5) n551 <= 1'b0; else if (1'b1) n551 <= n2095;
/* FF 18 12  5 */ always @(posedge n3, posedge n5) if (n5) n1174 <= 1'b0; else if (n1298) n1174 <= n2096;
/* FF 14 12  1 */ assign n553 = n2097;
/* FF 19 23  4 */ always @(posedge n3, posedge n5) if (n5) n1402 <= 1'b0; else if (1'b1) n1402 <= n2098;
/* FF 19 10  7 */ always @(posedge n3, posedge n5) if (n5) n951 <= 1'b0; else if (n580) n951 <= n2099;
/* FF 22 16  2 */ assign n1660 = n2100;
/* FF 26 17  2 */ always @(posedge n1, posedge n5) if (n5) n984 <= 1'b0; else if (n8) n984 <= n2101;
/* FF 14 19  5 */ always @(posedge n3, posedge n5) if (n5) n515 <= 1'b0; else if (1'b1) n515 <= n2102;
/* FF 17 14  1 */ assign n959 = n2103;
/* FF 19 24  2 */ always @(posedge n3, posedge n5) if (n5) n1407 <= 1'b0; else if (n1025) n1407 <= n2104;
/* FF 11 20  4 */ assign n391 = n2105;
/* FF 16 18  0 */ always @(posedge n3, posedge n5) if (n5) n979 <= 1'b0; else if (n800) n979 <= n2106;
/* FF 15 15  2 */ always @(posedge n3, posedge n5) if (n5) n787 <= 1'b0; else if (n944) n787 <= n2107;
/* FF 20 22  1 */ assign n2108 = n1618;
/* FF 10 19  1 */ always @(posedge n3, posedge n5) if (n5) n248 <= 1'b0; else if (n359) n248 <= n2109;
/* FF 13 11  0 */ assign n557 = n674;
/* FF 13 22  7 */ assign n639 = n2110;
/* FF 18 15  4 */ assign n2111 = n1334;
/* FF 14 15  0 */ assign n692 = n2112;
/* FF 19 11  4 */ always @(posedge n3, posedge n5) if (n5) n1178 <= 1'b0; else if (n1300) n1178 <= n2113;
/* FF 22 19  3 */ always @(posedge n3, posedge n5) if (n5) n1676 <= 1'b0; else if (n1369) n1676 <= n2114;
/* FF 17 15  6 */ assign n1090 = n2115;
/* FF 11 21  3 */ assign n273 = n2116;
/* FF 16 17  1 */ always @(posedge n3, posedge n5) if (n5) n974 <= 1'b0; else if (n702) n974 <= n2117;
/* FF 22 13  3 */ assign n2118 = n1714;
/* FF  6  8  1 */ assign io_28_0_0 = n2119;
/* FF 20 21  0 */ assign n1492 = n2120;
/* FF 16 15  0 */ assign n590 = n1097;
/* FF 23 13  4 */ assign n950 = n2121;
/* FF 24 14  4 */ always @(posedge n3, posedge n5) if (n5) n1590 <= 1'b0; else if (n467) n1590 <= n2122;
/* FF 13 12  1 */ assign n565 = n2123;
/* FF 14 21  6 */ always @(posedge n3, posedge n5) if (n5) n720 <= 1'b1; else if (n629) n720 <= n2124;
/* FF 12 20  0 */ always @(posedge n3, posedge n5) if (n5) n518 <= 1'b0; else if (n538) n518 <= n2125;
/* FF 17 11  3 */ assign n2126 = n1169;
/* FF 19 21  2 */ always @(posedge n3, posedge n5) if (n5) n1288 <= 1'b1; else if (n1145) n1288 <= n2127;
/* FF 23 14  6 */ always @(posedge n3, posedge n5) if (n5) n941 <= 1'b0; else if (n127) n941 <= n2128;
/* FF 24 17  2 */ always @(posedge n3, posedge n5) if (n5) n1360 <= 1'b0; else if (n1454) n1360 <= n2129;
/* FF 21 10  3 */ assign n1536 = n2130;
/* FF 12 10  1 */ assign n2131 = n555;
/* FF 11 18  2 */ assign n368 = n2132;
/* FF 22 12  0 */ always @(posedge n3, posedge n5) if (n5) n1632 <= 1'b0; else if (n1077) n1632 <= n2133;
/* FF 13 16  4 */ always @(posedge n3, posedge n5) if (n5) n586 <= 1'b0; else if (n492) n586 <= n2134;
/* FF 18 18  0 */ assign n1222 = n2135;
/* FF  6 11  0 */ always @(posedge n1, posedge n5) if (n5) n67 <= 1'b1; else if (1'b1) n67 <= n2136;
/* FF 23 18  0 */ always @(posedge n3, posedge n5) if (n5) n1733 <= 1'b0; else if (n1117) n1733 <= n2137;
/* FF 14 10  4 */ always @(posedge n1, posedge n5) if (n5) n662 <= 1'b0; else if (n672) n662 <= n2138;
/* FF 16 14  3 */ always @(posedge n3, posedge n5) if (n5) n943 <= 1'b0; else if (n321) n943 <= n2139;
/* FF  5 17  1 */ always @(posedge n3, posedge n5) if (n5) n46 <= 1'b0; else if (n4) n46 <= n2140;
/* FF 13 13  2 */ assign n320 = n2141;
/* FF 14 20  5 */ always @(posedge n3, posedge n5) if (n5) n396 <= 1'b0; else if (1'b1) n396 <= n2142;
/* FF 17 20  2 */ assign n1121 = n2143;
/* FF 19 18  3 */ assign n2144 = n1488;
/* FF 23 15  5 */ always @(posedge n3, posedge n5) if (n5) n1721 <= 1'b0; else if (n1654) n1721 <= n2145;
/* FF 21 16  5 */ assign n2146 = n1665;
/* FF 21 11  4 */ always @(posedge n3, posedge n5) if (n5) n1544 <= 1'b0; else if (n1631) n1544 <= n2147;
/* FF 18 22  5 */ always @(posedge n3, posedge n5) if (n5) n1259 <= 1'b0; else if (1'b1) n1259 <= n2148;
/* FF 17  9  4 */ always @(posedge n1, posedge n5) if (n5) n766 <= 1'b0; else if (n672) n766 <= n2149;
/* FF 11 19  1 */ assign n376 = n2150;
/* FF 10  9  1 */ always @(posedge n1, posedge n5) if (n5) n195 <= 1'b0; else if (1'b1) n195 <= n2151;
/* FF 22 15  1 */ assign n1652 = n2152;
/* FF 13 17  7 */ assign n594 = n2153;
/* FF 18 21  1 */ always @(posedge n3) if (n881) io_33_23_1 <= 1'b0 ? 1'b0 : n2154;
/* FF 19 14  6 */ assign n1318 = n2155;
/* FF 16 13  2 */ assign n935 = n2156;
/* FF  5 18  0 */ always @(posedge n3, posedge n5) if (n5) n52 <= 1'b0; else if (n4) n52 <= n2157;
/* FF 10 20  4 */ always @(posedge n3, posedge n5) if (n5) n263 <= 1'b0; else if (n144) n263 <= n2158;
/* FF 18  7  0 */ always @(posedge n3, posedge n5) if (n5) n654 <= 1'b0; else if (1'b1) n654 <= n2159;
/* FF 21 15  1 */ assign n2160 = n1657;
/* FF 20 25  1 */ always @(posedge n3, posedge n5) if (n5) n1415 <= 1'b0; else if (n1453) n1415 <= n2161;
/* FF 19 19  0 */ always @(posedge n3, posedge n5) if (n5) n969 <= 1'b0; else if (n985) n969 <= n2162;
/* FF 23 12  4 */ always @(posedge n3) if (n1301) n1491 <= 1'b0 ? 1'b0 : n2163;
/* FF 21 17  6 */ assign n1084 = n2164;
/* FF 21 12  5 */ always @(posedge n3, posedge n5) if (n5) n1550 <= 1'b0; else if (n1186) n1550 <= n2165;
/* FF 18 25  4 */ assign n1277 = n2166;
/* FF 17 10  5 */ always @(posedge n1, posedge n5) if (n5) n760 <= 1'b0; else if (n8) n760 <= n2167;
/* FF 11 16  0 */ assign n2168 = n489;
/* FF 22 14  6 */ always @(posedge n3, posedge n5) if (n5) n783 <= 1'b0; else if (n1651) n783 <= n2169;
/* FF 13 18  6 */ assign n512 = n2170;
/* FF 18 20  2 */ assign n1245 = n2171;
/* FF 23 16  2 */ always @(posedge n3, posedge n5) if (n5) n1152 <= 1'b0; else if (n1653) n1152 <= n2172;
/* FF 11 14  3 */ assign n315 = n2173;
/* FF 16  7  4 */ always @(negedge io_0_6_1, posedge n5) if (n5) n904 <= 1'b0; else if (1'b1) n904 <= n2174;
/* FF 19 15  5 */ always @(posedge n3, posedge n5) if (n5) n1329 <= 1'b0; else if (n619) n1329 <= n2175;
/* FF 16 12  5 */ always @(posedge n3, posedge n5) if (n5) n59 <= 1'b0; else if (n321) n59 <= n2176;
/* FF 15 26  2 */ always @(posedge n3, posedge n5) if (n5) n882 <= 1'b0; else if (n2) n882 <= n2177;
/* FF 12 12  4 */ always @(posedge io_0_6_1, posedge n5) if (n5) n427 <= 1'b0; else if (n563) n427 <= n2178;
/* FF 14 22  3 */ always @(posedge n3, posedge n5) if (n5) n724 <= 1'b0; else if (n704) n724 <= n2179;
/* FF 17 22  0 */ assign n1129 = n2180;
/* FF 19 16  1 */ always @(posedge n3, posedge n5) if (n5) n1321 <= 1'b0; else if (n949) n1321 <= n2182;
/* FF 22 10  3 */ always @(posedge n1, posedge n5) if (n5) n1624 <= 1'b0; else if (1'b1) n1624 <= n2183;
/* FF  7 11  6 */ always @(posedge n1, posedge n5) if (n5) n107 <= 1'b0; else if (1'b1) n107 <= n2184;
/* FF 21 18  7 */ assign n1596 = n2185;
/* FF 21 13  6 */ assign n1554 = n2186;
/* FF 12 15  6 */ assign n465 = n2187;
/* FF 18 24  7 */ assign n1241 = n2188;
/* FF 15  7  3 */ assign n736 = n907;
/* FF 13 19  1 */ assign n186 = n2189;
/* FF 15 21  0 */ assign n869 = n2190;
/* FF 18 23  3 */ always @(posedge n3) if (n881) io_33_5_1 <= 1'b0 ? 1'b0 : n2191;
/* FF 23 17  5 */ always @(posedge n3, posedge n5) if (n5) n1729 <= 1'b0; else if (n619) n1729 <= n2192;
/* FF 11 15  0 */ assign n323 = n2193;
/* FF 19 12  4 */ assign n1301 = n2194;
/* FF  9 19  2 */ assign io_0_30_0 = n2195;
/* FF 12 19  5 */ always @(posedge n3, posedge n5) if (n5) n508 <= 1'b1; else if (n620) n508 <= n2196;
/* FF 14 17  2 */ assign n708 = n2197;
/* FF 17 12  6 */ assign n1068 = n2198;
/* FF 17 23  7 */ assign n1144 = n2199;
/* FF 22 21  1 */ always @(posedge n3, posedge n5) if (n5) n1691 <= 1'b0; else if (n1652) n1691 <= n2200;
/* FF 21 19  0 */ assign n2201 = n1680;
/* FF 13 23  6 */ assign n2202 = n2203;
/* FF 21 14  7 */ assign n1562 = n2204;
/* FF  9 16  4 */ assign n169 = n2205;
/* FF 12 14  5 */ assign n447 = n2206;
/* FF 10 10  4 */ always @(posedge n1, posedge n5) if (n5) n200 <= 1'b0; else if (1'b1) n200 <= n2207;
/* FF 16 23  3 */ always @(posedge n3, posedge n5) if (n5) n1017 <= 1'b0; else if (n1010) n1017 <= n2208;
/* FF 10 17  6 */ assign n2209 = n2210;
/* FF 13 20  0 */ assign n621 = n2211;
/* FF 15 10  1 */ always @(posedge n1, posedge n5) if (n5) n748 <= 1'b0; else if (1'b1) n748 <= n2212;
/* FF 20 19  2 */ always @(posedge n3, posedge n5) if (n5) n1486 <= 1'b0; else if (n803) n1486 <= n2213;
/* FF 11 12  1 */ always @(posedge n3, posedge n5) if (n5) n212 <= 1'b0; else if (n26) n212 <= n2214;
/* FF 17 19  4 */ assign n2215 = n2216;
/* FF 19 13  3 */ assign n1304 = n2217;
/* FF 16 10  7 */ always @(posedge n1, posedge n5) if (n5) n668 <= 1'b0; else if (n672) n668 <= n2218;
/* FF 15 24  0 */ always @(posedge n3, posedge n5) if (n5) n886 <= 1'b0; else if (n2) n886 <= n2219;
/* FF 12 18  6 */ always @(posedge n3) if (1'b1) n500 <= n128 ? 1'b0 : n2220;
/* FF 17 13  5 */ assign n1075 = n2221;
/* FF 14 16  1 */ always @(posedge n3, posedge n5) if (n5) n698 <= 1'b0; else if (1'b1) n698 <= n2222;
/* FF 17 16  6 */ assign n713 = n2223;
/* FF 22 20  2 */ assign n2224 = n1740;
/* FF 10 14  1 */ always @(posedge n1) if (1'b1) n213 <= n7 ? 1'b0 : n2225;
/* FF 21 20  1 */ always @(posedge n3, posedge n5) if (n5) n1603 <= 1'b0; else if (n270) n1603 <= n2226;
/* FF 13 24  7 */ assign n2227 = n2228;
/* FF  9 17  7 */ always @(posedge n3, posedge n5) if (n5) n175 <= 1'b1; else if (n172) n175 <= n2229;
/* FF 12 13  4 */ always @(posedge n3, posedge n5) if (n5) n435 <= 1'b0; else if (n573) n435 <= n2230;
/* FF 20 12  0 */ always @(posedge n3, posedge n5) if (n5) n1431 <= 1'b0; else if (n1299) n1431 <= n2231;
/* FF 10 13  5 */ always @(posedge n1, posedge n5) if (n5) n209 <= 1'b0; else if (n138) n209 <= n2232;
/* FF 16 22  0 */ always @(posedge n3) if (n881) io_33_30_0 <= 1'b0 ? 1'b0 : n2233;
/* FF 10 16  5 */ always @(posedge n1) if (1'b1) n235 <= n7 ? 1'b0 : n2234;
/* FF 13 21  3 */ assign n257 = n2235;
/* FF 20 18  1 */ always @(posedge n3, posedge n5) if (n5) n1480 <= 1'b0; else if (n1369) n1480 <= n2236;
/* FF 11 13  6 */ always @(posedge n3, posedge n5) if (n5) n303 <= 1'b0; else if (n441) n303 <= n2237;
/* FF 19 10  2 */ always @(posedge n3, posedge n5) if (n5) n1290 <= 1'b0; else if (n580) n1290 <= n2238;
/* FF 15 25  7 */ always @(posedge n3, posedge n5) if (n5) n897 <= 1'b0; else if (n2) n897 <= n2239;
/* FF  7 13  5 */ always @(posedge n1, posedge n5) if (n5) n124 <= 1'b0; else if (1'b1) n124 <= n2240;
/* FF 12 17  7 */ always @(posedge n3) if (1'b1) n491 <= n128 ? 1'b0 : n2241;
/* FF 14 19  0 */ always @(posedge n3, posedge n5) if (n5) n269 <= 1'b0; else if (1'b1) n269 <= n2242;
/* FF 17 14  4 */ assign n1081 = n2243;
/* FF 17 17  5 */ assign n2244 = n1221;
/* FF 22 23  3 */ always @(posedge n3, posedge n5) if (n5) n1694 <= 1'b0; else if (n1656) n1694 <= n2245;
/* FF 21 21  2 */ assign n1566 = n2246;
/* FF 11  9  3 */ assign n276 = n407;
/* FF 16 21  1 */ always @(posedge n3, posedge n5) if (n5) n999 <= 1'b0; else if (n995) n999 <= n2247;
/* FF 10 19  4 */ always @(posedge n3, posedge n5) if (n5) n251 <= 1'b0; else if (n359) n251 <= n2248;
/* FF 13 22  2 */ assign n634 = n2249;
/* FF  6 12  1 */ assign n76 = n2250;
/* FF 20 17  0 */ assign n1094 = n2251;
/* FF 23 20  6 */ always @(posedge n3, posedge n5) if (n5) n1505 <= 1'b0; else if (n1655) n1505 <= n2252;
/* FF 11 10  7 */ always @(posedge n1, posedge n5) if (n5) n285 <= 1'b1; else if (1'b1) n285 <= n2253;
/* FF 19 11  1 */ always @(posedge n3, posedge n5) if (n5) n1295 <= 1'b0; else if (n1300) n1295 <= n2254;
/* FF 12 16  0 */ assign n481 = n2255;
/* FF 17 15  3 */ assign n2256 = n1206;
/* FF 19 25  2 */ always @(posedge n3, posedge n5) if (n5) n1411 <= 1'b0; else if (n1012) n1411 <= n2257;
/* FF 17 18  4 */ assign n2258 = n2259;
/* FF 22 13  6 */ assign n2260 = n1715;
/* FF  7 15  2 */ always @(posedge n1, posedge n5) if (n5) io_0_27_1 <= 1'b0; else if (1'b1) io_0_27_1 <= n2261;
/* FF 21 22  3 */ assign n1610 = n2262;
/* FF 11 22  2 */ always @(posedge n3, posedge n5) if (n5) n400 <= 1'b1; else if (n273) n400 <= n2263;
/* FF 16 15  7 */ assign n688 = n2264;
/* FF 10 15  7 */ always @(posedge n1) if (1'b1) n226 <= n7 ? 1'b0 : n2265;
/* FF 16 20  6 */ assign n144 = n2266;
/* FF 15 18  5 */ always @(posedge n3, posedge n5) if (n5) n822 <= 1'b0; else if (n826) n822 <= n2267;
/* FF 18 14  0 */ assign n2268 = n1324;
/* FF 20 16  7 */ always @(posedge n3, posedge n5) if (n5) n1211 <= 1'b0; else if (n1455) n1211 <= n2269;
/* FF 12 20  5 */ always @(posedge n3, posedge n5) if (n5) n521 <= 1'b0; else if (n538) n521 <= n2270;
/* FF 11 11  4 */ always @(posedge n1, posedge n5) if (n5) n280 <= 1'b0; else if (1'b1) n280 <= n2271;
/* FF 22 18  1 */ assign n2272 = n1737;
/* FF 13  9  2 */ always @(posedge n3, posedge n5) if (n5) n547 <= 1'b0; else if (1'b1) n547 <= n2273;
/* FF 21 10  6 */ always @(posedge n1, posedge n5) if (n5) n1538 <= 1'b0; else if (1'b1) n1538 <= n2274;
/* FF 12 23  1 */ assign n2275 = n2276;
/* FF 17  8  2 */ always @(posedge n3, posedge n5) if (n5) n747 <= 1'b0; else if (1'b1) n747 <= n2277;
/* FF 19 22  3 */ always @(posedge n3, posedge n5) if (n5) n1392 <= 1'b0; else if (1'b1) n1392 <= n2278;
/* FF 22 17  5 */ assign n1668 = n2279;
/* FF 16 16  3 */ always @(posedge n3, posedge n5) if (n5) n964 <= 1'b0; else if (n799) n964 <= n2280;
/* FF 22 12  5 */ always @(posedge n3, posedge n5) if (n5) n1637 <= 1'b0; else if (n1077) n1637 <= n2281;
/* FF 15 13  1 */ assign n775 = n946;
/* FF 20 20  4 */ always @(posedge n3, posedge n5) if (n5) n1384 <= 1'b0; else if (n996) n1384 <= n2282;
/* FF 16 14  4 */ assign n609 = n2283;
/* FF 16 19  7 */ always @(posedge n3, posedge n5) if (n5) n992 <= 1'b1; else if (n801) n992 <= n2284;
/* FF 15 19  6 */ always @(posedge n3, posedge n5) if (n5) n841 <= 1'b0; else if (n629) n841 <= n2285;
/* FF 15 14  5 */ always @(posedge n3, posedge n5) if (n5) n771 <= 1'b0; else if (1'b1) n771 <= n2286;
/* FF 18 17  1 */ assign n2287 = n1352;
/* FF 20 23  6 */ always @(posedge n3) if (n688) n1521 <= 1'b0 ? 1'b0 : n2288;
/* FF 24 16  2 */ always @(posedge n3, posedge n5) if (n5) n1210 <= 1'b0; else if (n619) n1210 <= n2289;
/* FF 21 11  1 */ always @(posedge n3, posedge n5) if (n5) n1541 <= 1'b0; else if (n1631) n1541 <= n2290;
/* FF 12 22  2 */ assign n2291 = n2292;
/* FF 19 23  0 */ always @(posedge n3, posedge n5) if (n5) n1024 <= 1'b0; else if (1'b1) n1024 <= n2293;
/* FF 22 16  6 */ assign n2294 = n1725;
/* FF 22 15  4 */ assign n1631 = n2295;
/* FF 20 11  5 */ always @(posedge n3, posedge n5) if (n5) n1095 <= 1'b0; else if (n1199) n1095 <= n2296;
/* FF 19 24  6 */ always @(posedge n3, posedge n5) if (n5) n796 <= 1'b0; else if (n1025) n796 <= n2297;
/* FF 11 20  0 */ assign n387 = n2298;
/* FF 16 13  5 */ assign n596 = n2299;
/* FF 16 18  4 */ always @(posedge n3, posedge n5) if (n5) n982 <= 1'b0; else if (n800) n982 <= n2300;
/* FF 10 20  1 */ always @(posedge n3, posedge n5) if (n5) n260 <= 1'b0; else if (n144) n260 <= n2301;
/* FF 15 16  7 */ assign n801 = n2302;
/* FF 21 15  6 */ assign n1575 = n2303;
/* FF 15 15  6 */ always @(posedge n3, posedge n5) if (n5) n790 <= 1'b0; else if (n944) n790 <= n2304;
/* FF 18 16  2 */ always @(posedge n1, posedge n5) if (n5) n595 <= 1'b0; else if (n8) n595 <= n2305;
/* FF  6  9  6 */ assign n64 = n2306;
/* FF 20 22  5 */ always @(posedge n3, posedge n5) if (n5) n1273 <= 1'b0; else if (1'b1) n1273 <= n2307;
/* FF 17 24  1 */ assign n2308 = n2309;
/* FF 24 15  3 */ always @(posedge n3, posedge n5) if (n5) n1204 <= 1'b0; else if (n958) n1204 <= n2310;
/* FF 13 11  4 */ assign n561 = n675;
/* FF 21 12  0 */ always @(posedge n3, posedge n5) if (n5) n1545 <= 1'b0; else if (n1186) n1545 <= n2311;
/* FF 12 21  3 */ assign n533 = n2312;
/* FF 17 10  0 */ always @(posedge n1, posedge n5) if (n5) n930 <= 1'b0; else if (n8) n930 <= n2313;
/* FF 19 20  1 */ always @(posedge n3, posedge n5) if (n5) n1377 <= 1'b0; else if (1'b1) n1377 <= n2314;
/* FF 22 19  7 */ assign n1678 = n2315;
/* FF 22 14  3 */ always @(posedge n3, posedge n5) if (n5) n1647 <= 1'b0; else if (n1651) n1647 <= n2316;
/* FF 23 16  5 */ always @(posedge n3, posedge n5) if (n5) n1598 <= 1'b0; else if (n1653) n1598 <= n2317;
/* FF 11 14  6 */ assign n318 = n2318;
/* FF 16 12  2 */ assign n2319 = n1070;
/* FF 16 17  5 */ always @(posedge n3, posedge n5) if (n5) n975 <= 1'b0; else if (n702) n975 <= n2320;
/* FF 13 15  1 */ always @(posedge n3) if (io_0_25_1) n578 <= 1'b0 ? 1'b0 : n2321;
/* FF 15 17  0 */ always @(posedge n3, posedge n5) if (n5) n808 <= 1'b0; else if (n609) n808 <= n2322;
/* FF 15 12  7 */ always @(posedge n3, posedge n5) if (n5) n14 <= 1'b0; else if (1'b1) n14 <= n2323;
/* FF 18 19  3 */ assign n1234 = n2324;
/* FF 20 21  4 */ assign n1112 = n2325;
/* FF 24 14  0 */ always @(posedge n3, posedge n5) if (n5) n1104 <= 1'b0; else if (n467) n1104 <= n2326;
/* FF 13 12  5 */ always @(posedge io_0_6_1, posedge n5) if (n5) n569 <= 1'b0; else if (1'b1) n569 <= n2327;
/* FF 21 13  3 */ assign n1552 = n2328;
/* FF 19 21  6 */ always @(posedge n3, posedge n5) if (n5) n1285 <= 1'b0; else if (n1145) n1285 <= n2329;
/* FF 11 17  4 */ assign n355 = n497;
/* FF 24 17  6 */ always @(posedge n3, posedge n5) if (n5) n1742 <= 1'b0; else if (n1454) n1742 <= n2330;
/* FF 15 21  5 */ assign n874 = n2331;
/* FF 20  9  7 */ assign n1424 = n2332;
/* FF 23 17  2 */ assign n1727 = n2333;
/* FF 11 15  5 */ assign n328 = n2334;
/* FF 11 18  6 */ assign n372 = n2335;
/* FF 16 11  3 */ always @(posedge n3, posedge n5) if (n5) n202 <= 1'b0; else if (n938) n202 <= n2336;
/* FF 13 16  0 */ always @(posedge n3, posedge n5) if (n5) n582 <= 1'b0; else if (n492) n582 <= n2337;
/* FF 15 22  1 */ assign n2338 = n2339;
/* FF 18  9  5 */ always @(posedge n3, posedge n5) if (n5) n1156 <= 1'b0; else if (n215) n1156 <= n2340;
/* FF 18 18  4 */ assign n1225 = n2341;
/* FF  6 11  4 */ always @(posedge n1, posedge n5) if (n5) n71 <= 1'b0; else if (1'b1) n71 <= n2342;
/* FF 14 10  0 */ always @(posedge n1, posedge n5) if (n5) n658 <= 1'b0; else if (n672) n658 <= n2343;
/* FF 19 17  3 */ assign n1346 = n2344;
/* FF 22 21  4 */ always @(posedge n3, posedge n5) if (n5) n1383 <= 1'b0; else if (n1652) n1383 <= n2345;
/* FF 24 13  1 */ always @(posedge n3, posedge n5) if (n5) n1712 <= 1'b0; else if (n805) n1712 <= n2346;
/* FF 13 13  6 */ always @(posedge io_0_6_1, posedge n5) if (n5) n36 <= 1'b0; else if (n563) n36 <= n2347;
/* FF 21 14  2 */ always @(posedge n3, posedge n5) if (n5) n1559 <= 1'b0; else if (n805) n1559 <= n2348;
/* FF  9 16  3 */ assign n168 = n2349;
/* FF 14 20  1 */ always @(posedge n3, posedge n5) if (n5) n397 <= 1'b0; else if (1'b1) n397 <= n2350;
/* FF 19 18  7 */ assign n1359 = n2351;
/* FF 10 10  1 */ assign n197 = n2352;
/* FF 16 23  6 */ always @(posedge n3, posedge n5) if (n5) n1020 <= 1'b0; else if (n1010) n1020 <= n2353;
/* FF 21 16  1 */ assign n2354 = n1663;
/* FF 15 10  4 */ always @(posedge n1, posedge n5) if (n5) n753 <= 1'b0; else if (1'b1) n753 <= n2355;
/* FF 11 12  4 */ always @(posedge n3, posedge n5) if (n5) n35 <= 1'b0; else if (n26) n35 <= n2356;
/* FF 11 19  5 */ assign n380 = n2357;
/* FF 16 10  0 */ always @(posedge n1, posedge n5) if (n5) n918 <= 1'b0; else if (n672) n918 <= n2358;
/* FF  9 12  5 */ assign n156 = n2359;
/* FF 13 17  3 */ assign n374 = n711;
/* FF 18 21  5 */ always @(posedge n3) if (n881) io_26_33_0 <= 1'b0 ? 1'b0 : n2360;
/* FF 19 14  2 */ assign n1317 = n2361;
/* FF 22 20  7 */ assign n1688 = n2362;
/* FF 16 24  4 */ always @(posedge n3, posedge n5) if (n5) n192 <= 1'b0; else if (n1010) n192 <= n2363;
/* FF  9 17  0 */ assign n172 = n2364;
/* FF 20 12  5 */ always @(posedge n3, posedge n5) if (n5) n1309 <= 1'b0; else if (n1299) n1309 <= n2365;
/* FF 19 19  4 */ always @(posedge n3, posedge n5) if (n5) n961 <= 1'b0; else if (n985) n961 <= n2366;
/* FF 10 13  0 */ always @(posedge n1, posedge n5) if (n5) n203 <= 1'b0; else if (n138) n203 <= n2367;
/* FF 16 22  5 */ assign n5 = n2368;
/* FF 22 11  0 */ always @(posedge n1, posedge n5) if (n5) n1627 <= 1'b0; else if (1'b1) n1627 <= n2369;
/* FF 21 17  2 */ assign n1586 = n2370;
/* FF 20 15  1 */ assign n1454 = n2371;
/* FF 11 13  3 */ always @(posedge n3, posedge n5) if (n5) n300 <= 1'b0; else if (n441) n300 <= n2372;
/* FF 11 16  4 */ assign n341 = n2373;
/* FF 16  9  1 */ always @(posedge n3, posedge n5) if (n5) n756 <= 1'b0; else if (n933) n756 <= n2374;
/* FF 13 18  2 */ assign n142 = n2375;
/* FF 15 20  3 */ assign n856 = n2376;
/* FF 18 20  6 */ always @(posedge n3, posedge n5) if (n5) n1248 <= 1'b0; else if (n704) n1248 <= n2377;
/* FF 16  7  0 */ always @(negedge io_0_6_1, posedge n5) if (n5) n900 <= 1'b0; else if (1'b1) n900 <= n2378;
/* FF 19 15  1 */ assign n2380 = n1463;
/* FF 22 23  6 */ always @(posedge n3, posedge n5) if (n5) n1361 <= 1'b0; else if (n1656) n1361 <= n2381;
/* FF 24 22  4 */ assign io_33_27_1 = n2382;
/* FF  9 18  1 */ always @(posedge n3, posedge n5) if (n5) n177 <= 1'b0; else if (n172) n177 <= n2383;
/* FF 12 12  0 */ always @(posedge io_0_6_1, posedge n5) if (n5) n423 <= 1'b0; else if (n563) n423 <= n2384;
/* FF 19 16  5 */ always @(posedge n3, posedge n5) if (n5) n1338 <= 1'b0; else if (n949) n1338 <= n2385;
/* FF 16 21  4 */ always @(posedge n3, posedge n5) if (n5) n1002 <= 1'b0; else if (n995) n1002 <= n2386;
/* FF 16 26  5 */ always @(posedge n3, posedge n5) if (n5) n1044 <= 1'b0; else if (n704) n1044 <= n2387;
/* FF 21 18  3 */ assign n2388 = n1674;
/* FF 15  7  7 */ always @(negedge io_0_6_1, posedge n5) if (n5) n740 <= 1'b0; else if (1'b1) n740 <= n2389;
/* FF 18 24  3 */ assign n2390 = n1413;
/* FF 20 14  2 */ always @(posedge n1, posedge n5) if (n5) n1055 <= 1'b0; else if (n8) n1055 <= n2391;
/* FF 23 20  1 */ always @(posedge n3, posedge n5) if (n5) n1229 <= 1'b0; else if (n1655) n1229 <= n2392;
/* FF 11 10  2 */ assign n2393 = n413;
/* FF  9 14  7 */ assign n80 = n2394;
/* FF 13 19  5 */ assign n618 = n2395;
/* FF 18 23  7 */ always @(posedge n3) if (n881) io_33_21_0 <= 1'b0 ? 1'b0 : n2396;
/* FF 14 18  4 */ always @(posedge n3, posedge n5) if (n5) n183 <= 1'b0; else if (1'b1) n183 <= n2397;
/* FF 14  7  3 */ always @(negedge io_0_6_1, posedge n5) if (n5) n649 <= 1'b0; else if (1'b1) n649 <= n2398;
/* FF 19 12  0 */ assign n1186 = n2399;
/* FF 22 22  1 */ always @(posedge n3, posedge n5) if (n5) n1697 <= 1'b0; else if (n1010) n1697 <= n2400;
/* FF 12 19  1 */ always @(posedge n3, posedge n5) if (n5) n504 <= 1'b0; else if (n620) n504 <= n2401;
/* FF 17 12  2 */ assign n1064 = n2402;
/* FF 10 15  2 */ always @(posedge n1) if (1'b1) n221 <= n7 ? 1'b0 : n2403;
/* FF 16 20  3 */ assign n270 = n2404;
/* FF 21 19  4 */ assign n2405 = n1683;
/* FF 13 23  2 */ assign n2406 = n2407;
/* FF 15  9  1 */ always @(posedge n3, posedge n5) if (n5) n653 <= 1'b0; else if (1'b1) n653 <= n2408;
/* FF 18 14  5 */ assign n1192 = n2409;
/* FF 20 13  3 */ assign n2410 = n1558;
/* FF 11 11  1 */ assign n293 = n2411;
/* FF 22 18  6 */ assign n1671 = n2412;
/* FF 10 17  2 */ always @(posedge n1) if (1'b1) n241 <= n7 ? 1'b0 : n2413;
/* FF  9 15  0 */ assign n160 = n2414;
/* FF 13 20  4 */ assign n625 = n2415;
/* FF 18 13  1 */ always @(posedge n1, posedge n5) if (n5) n758 <= 1'b0; else if (n8) n758 <= n2416;
/* FF 14 13  5 */ always @(posedge n3, posedge n5) if (n5) n687 <= 1'b0; else if (n690) n687 <= n2417;
/* FF 19 22  6 */ always @(posedge n3, posedge n5) if (n5) n1395 <= 1'b0; else if (1'b1) n1395 <= n2418;
/* FF 17 19  0 */ assign n2419 = n2420;
/* FF 19 13  7 */ assign n1307 = n2421;
/* FF 22 17  0 */ assign n2422 = n1730;
/* FF 15 13  6 */ always @(posedge n3, posedge n5) if (n5) n778 <= 1'b0; else if (n321) n778 <= n2423;
/* FF 12 18  2 */ always @(posedge n3) if (1'b1) n486 <= n128 ? 1'b0 : n2424;
/* FF 14 16  5 */ always @(posedge n3, posedge n5) if (n5) n322 <= 1'b1; else if (1'b1) n322 <= n2425;
/* FF 17 13  1 */ assign n2426 = n1187;
/* FF 16 19  2 */ always @(posedge n3, posedge n5) if (n5) n877 <= 1'b1; else if (n801) n877 <= n2427;
/* FF 21 20  5 */ always @(posedge n3, posedge n5) if (n5) n1606 <= 1'b0; else if (n270) n1606 <= n2428;
/* FF 13 24  3 */ assign n2429 = n2430;
/* FF 15 14  0 */ assign n769 = n955;
/* FF 18 17  4 */ assign n2431 = n1353;
/* FF 18 26  5 */ assign n1280 = n2432;
/* FF 10 16  1 */ always @(posedge n1) if (1'b1) n231 <= n7 ? 1'b0 : n2433;
/* FF 13 21  7 */ assign n630 = n2434;
/* FF 18 12  2 */ always @(posedge n3, posedge n5) if (n5) n1165 <= 1'b0; else if (n1298) n1165 <= n2435;
/* FF 14 12  6 */ always @(posedge n3) if (1'b1) n28 <= 1'b0 ? 1'b0 : n2436;
/* FF 19 23  5 */ always @(posedge n3, posedge n5) if (n5) n1403 <= 1'b0; else if (1'b1) n1403 <= n2437;
/* FF 19 10  6 */ always @(posedge n3, posedge n5) if (n5) n954 <= 1'b0; else if (n580) n954 <= n2438;
/* FF 22 16  3 */ assign n2439 = n1723;
/* FF 12 17  3 */ always @(posedge n3) if (1'b1) n471 <= n128 ? 1'b0 : n2440;
/* FF 14 19  4 */ always @(posedge n3, posedge n5) if (n5) n187 <= 1'b0; else if (1'b1) n187 <= n2441;
/* FF 17 14  0 */ assign n2442 = n1196;
/* FF 19 24  1 */ always @(posedge n3, posedge n5) if (n5) n1406 <= 1'b0; else if (n1025) n1406 <= n2443;
/* FF 16 18  1 */ always @(posedge n3, posedge n5) if (n5) n843 <= 1'b0; else if (n800) n843 <= n2444;
/* FF 21 21  6 */ always @(posedge n3, posedge n5) if (n5) n1613 <= 1'b0; else if (n704) n1613 <= n2445;
/* FF 13 25  0 */ assign io_0_22_1 = n2446;
/* FF 15 15  3 */ always @(posedge n3, posedge n5) if (n5) n785 <= 1'b0; else if (n944) n785 <= n2447;
/* FF 10 19  0 */ always @(posedge n3, posedge n5) if (n5) n247 <= 1'b1; else if (n359) n247 <= n2448;
/* FF 13 11  1 */ assign n558 = n2449;
/* FF 13 22  6 */ assign n638 = n2450;
/* FF 18 15  3 */ assign n1201 = n2451;
/* FF 14 15  7 */ assign n691 = n2452;
/* FF 19 20  4 */ always @(posedge n3, posedge n5) if (n5) n1380 <= 1'b0; else if (1'b1) n1380 <= n2453;
/* FF 19 11  5 */ always @(posedge n3, posedge n5) if (n5) n1167 <= 1'b0; else if (n1300) n1167 <= n2454;
/* FF 22 19  2 */ assign n1348 = n2455;
/* FF 17 15  7 */ assign n1091 = n2456;
/* FF 16 17  0 */ always @(posedge n3, posedge n5) if (n5) n973 <= 1'b0; else if (n702) n973 <= n2457;
/* FF 22 13  2 */ always @(posedge n3, posedge n5) if (n5) n1639 <= 1'b0; else if (n805) n1639 <= n2458;
/* FF 15 12  2 */ assign n767 = n2459;
/* FF 18 19  6 */ assign n1237 = n2460;
/* FF 16 15  3 */ assign n238 = n1098;
/* FF 23 13  5 */ always @(posedge n3, posedge n5) if (n5) n1711 <= 1'b0; else if (n793) n1711 <= n2461;
/* FF 24 14  5 */ always @(posedge n3, posedge n5) if (n5) n1370 <= 1'b0; else if (n467) n1370 <= n2462;
/* FF  9 10  3 */ assign n150 = n2463;
/* FF 13 12  0 */ assign n2464 = n2465;
/* FF 15 18  1 */ always @(posedge n3, posedge n5) if (n5) n716 <= 1'b0; else if (n826) n716 <= n2467;
/* FF 14 14  0 */ always @(posedge n3, posedge n5) if (n5) n689 <= 1'b0; else if (n321) n689 <= n2468;
/* FF 17 11  4 */ assign n1059 = n2469;
/* FF 19 21  3 */ always @(posedge n3, posedge n5) if (n5) n1284 <= 1'b0; else if (n1145) n1284 <= n2470;
/* FF 23 14  1 */ always @(posedge n3, posedge n5) if (n5) n1462 <= 1'b0; else if (n127) n1462 <= n2471;
/* FF 24 17  1 */ always @(posedge n3, posedge n5) if (n5) n1483 <= 1'b0; else if (n1454) n1483 <= n2472;
/* FF 21 10  2 */ always @(posedge n1, posedge n5) if (n5) n1535 <= 1'b0; else if (1'b1) n1535 <= n2473;
/* FF 12 23  5 */ assign n2474 = n2475;
/* FF 22 12  1 */ always @(posedge n3, posedge n5) if (n5) n1633 <= 1'b0; else if (n1077) n1633 <= n2476;
/* FF 13 16  7 */ always @(posedge n3, posedge n5) if (n5) n589 <= 1'b0; else if (n492) n589 <= n2477;
/* FF  7 12  7 */ assign n122 = n2478;
/* FF 18 18  1 */ assign n2479 = n1363;
/* FF 20 20  0 */ always @(posedge n3, posedge n5) if (n5) n1114 <= 1'b0; else if (n996) n1114 <= n2480;
/* FF 23 18  3 */ always @(posedge n3, posedge n5) if (n5) n1250 <= 1'b0; else if (n1117) n1250 <= n2481;
/* FF 14 10  5 */ always @(posedge n1, posedge n5) if (n5) n663 <= 1'b0; else if (n672) n663 <= n2482;
/* FF 16 14  0 */ assign n704 = n2483;
/* FF  5 17  6 */ always @(posedge n3, posedge n5) if (n5) n50 <= 1'b0; else if (n4) n50 <= n2484;
/* FF 13 13  3 */ assign n572 = n2485;
/* FF 17 20  5 */ assign n1124 = n2486;
/* FF 19 18  2 */ assign n1356 = n2487;
/* FF 23 15  2 */ always @(posedge n3, posedge n5) if (n5) n1208 <= 1'b0; else if (n1654) n1208 <= n2488;
/* FF 21 16  4 */ assign n1581 = n2489;
/* FF 21 11  5 */ always @(posedge n3, posedge n5) if (n5) n570 <= 1'b0; else if (n1631) n570 <= n2490;
/* FF 18 22  6 */ always @(posedge n3, posedge n5) if (n5) n1260 <= 1'b0; else if (1'b1) n1260 <= n2491;
/* FF 12 22  6 */ assign n2492 = n2493;
/* FF 10  9  0 */ always @(posedge n1, posedge n5) if (n5) n194 <= 1'b0; else if (1'b1) n194 <= n2494;
/* FF 22 15  0 */ assign n1651 = n2495;
/* FF 13 17  4 */ assign n493 = n2496;
/* FF 18 21  0 */ always @(posedge n3) if (n881) io_33_21_1 <= 1'b0 ? 1'b0 : n2497;
/* FF 20 11  1 */ always @(posedge n3, posedge n5) if (n5) n1428 <= 1'b0; else if (n1199) n1428 <= n2498;
/* FF 16 13  1 */ always @(posedge n3, posedge n5) if (n5) n180 <= 1'b0; else if (n321) n180 <= n2499;
/* FF  5 18  7 */ always @(posedge n3, posedge n5) if (n5) n29 <= 1'b0; else if (n4) n29 <= n2500;
/* FF 10 20  5 */ always @(posedge n3, posedge n5) if (n5) n264 <= 1'b1; else if (n144) n264 <= n2501;
/* FF 15 16  3 */ assign n620 = n2502;
/* FF 21 15  2 */ assign n1572 = n2503;
/* FF 20 25  0 */ always @(posedge n3, posedge n5) if (n5) n1113 <= 1'b0; else if (n1453) n1113 <= n2504;
/* FF 17 21  6 */ assign n993 = n2505;
/* FF 19 19  1 */ always @(posedge n3, posedge n5) if (n5) n1366 <= 1'b0; else if (n985) n1366 <= n2506;
/* FF 17 24  5 */ assign n2507 = n2508;
/* FF 23 12  3 */ always @(posedge n3) if (n1301) n1709 <= 1'b0 ? 1'b0 : n2509;
/* FF 21 17  7 */ always @(posedge n3, posedge n5) if (n5) n1589 <= 1'b0; else if (n1179) n1589 <= n2510;
/* FF 21 12  4 */ always @(posedge n3, posedge n5) if (n5) n1549 <= 1'b0; else if (n1186) n1549 <= n2511;
/* FF 12 21  7 */ assign n537 = n2512;
/* FF 17 10  4 */ always @(posedge n1, posedge n5) if (n5) n757 <= 1'b0; else if (n8) n757 <= n2513;
/* FF 22 14  7 */ always @(posedge n3, posedge n5) if (n5) n784 <= 1'b0; else if (n1651) n784 <= n2514;
/* FF 13 18  5 */ assign n606 = n2515;
/* FF 23 16  1 */ always @(posedge n3, posedge n5) if (n5) n939 <= 1'b0; else if (n1653) n939 <= n2516;
/* FF 11 14  2 */ assign n314 = n2517;
/* FF 16 12  6 */ assign n932 = n1072;
/* FF  5 19  0 */ always @(posedge n3, posedge n5) if (n5) n60 <= 1'b0; else if (n4) n60 <= n2518;
/* FF 22 24  0 */ always @(posedge n3, posedge n5) if (n5) n1698 <= 1'b0; else if (n1369) n1698 <= n2519;
/* FF 15 17  4 */ always @(posedge n3, posedge n5) if (n5) n812 <= 1'b0; else if (n609) n812 <= n2520;
/* FF 20 24  7 */ assign n1524 = n2521;
/* FF 17 22  7 */ assign n1136 = n2522;
/* FF 14 11  3 */ always @(posedge n1, posedge n5) if (n5) n670 <= 1'b0; else if (1'b1) n670 <= n2523;
/* FF 19 16  0 */ always @(posedge n3, posedge n5) if (n5) n1332 <= 1'b0; else if (n949) n1332 <= n2524;
/* FF 22 10  4 */ always @(posedge n1, posedge n5) if (n5) n1294 <= 1'b0; else if (1'b1) n1294 <= n2525;
/* FF 21 18  6 */ assign n2526 = n1675;
/* FF 21 13  7 */ assign n1555 = n2527;
/* FF 12 15  1 */ assign n460 = n2528;
/* FF 15  7  0 */ assign n733 = n2529;
/* FF 18 24  4 */ assign n2530 = n1414;
/* FF 13 19  2 */ assign n143 = n2531;
/* FF 15 21  1 */ assign n870 = n2532;
/* FF 18 23  2 */ always @(posedge n3) if (n881) io_33_6_0 <= 1'b0 ? 1'b0 : n2533;
/* FF 23 17  6 */ assign n2534 = n1747;
/* FF 11 15  1 */ assign n324 = n2535;
/* FF 16 11  7 */ always @(posedge n3, posedge n5) if (n5) n928 <= 1'b0; else if (n938) n928 <= n2536;
/* FF  5 20  1 */ assign n7 = n2537;
/* FF 15 22  5 */ assign n2538 = n2539;
/* FF 18  9  1 */ always @(posedge n3, posedge n5) if (n5) n1157 <= 1'b0; else if (n215) n1157 <= n2540;
/* FF 12 19  4 */ always @(posedge n3, posedge n5) if (n5) n507 <= 1'b0; else if (n620) n507 <= n2541;
/* FF 17 23  0 */ assign n1137 = n2542;
/* FF 22 21  0 */ always @(posedge n3, posedge n5) if (n5) n1689 <= 1'b0; else if (n1652) n1689 <= n2543;
/* FF 21 19  1 */ assign n2544 = n1681;
/* FF 13 23  7 */ assign n2545 = n2546;
/* FF 21 14  6 */ assign n2547 = n1650;
/* FF  9 16  7 */ assign n170 = n2548;
/* FF 12 14  2 */ assign n444 = n2549;
/* FF 10 10  5 */ assign n2550 = n2551;
/* FF 16 23  2 */ always @(posedge n3, posedge n5) if (n5) n1016 <= 1'b0; else if (n1010) n1016 <= n2552;
/* FF 13 20  3 */ assign n624 = n2553;
/* FF 15 10  0 */ always @(posedge n1, posedge n5) if (n5) n752 <= 1'b0; else if (1'b1) n752 <= n2554;
/* FF 20 19  5 */ always @(posedge n3, posedge n5) if (n5) n1116 <= 1'b0; else if (n803) n1116 <= n2555;
/* FF 11 12  0 */ always @(posedge n3, posedge n5) if (n5) n159 <= 1'b0; else if (n26) n159 <= n2556;
/* FF 17 19  5 */ assign n2557 = n2558;
/* FF 16 10  4 */ always @(posedge n1, posedge n5) if (n5) n921 <= 1'b0; else if (n672) n921 <= n2559;
/* FF  9 12  1 */ always @(posedge n1, posedge n5) if (n5) n154 <= 1'b0; else if (1'b1) n154 <= n2560;
/* FF 15 24  7 */ always @(posedge n3, posedge n5) if (n5) n891 <= 1'b0; else if (n2) n891 <= n2561;
/* FF 12 18  7 */ always @(posedge n3) if (1'b1) n501 <= n128 ? 1'b0 : n2562;
/* FF 17 16  1 */ assign n1101 = n2563;
/* FF 22 20  3 */ assign n2564 = n1741;
/* FF 10 14  2 */ always @(posedge n1) if (1'b1) n214 <= n7 ? 1'b0 : n2565;
/* FF 16 24  0 */ always @(posedge n3, posedge n5) if (n5) n1022 <= 1'b0; else if (n1010) n1022 <= n2566;
/* FF 21 20  0 */ always @(posedge n3, posedge n5) if (n5) n1599 <= 1'b0; else if (n270) n1599 <= n2567;
/* FF 13 24  6 */ assign n2568 = n2569;
/* FF 12 13  3 */ always @(posedge n3, posedge n5) if (n5) n434 <= 1'b1; else if (n573) n434 <= n2570;
/* FF 20 12  1 */ always @(posedge n3, posedge n5) if (n5) n1432 <= 1'b0; else if (n1299) n1432 <= n2571;
/* FF 10 13  4 */ always @(posedge n1, posedge n5) if (n5) n204 <= 1'b0; else if (n138) n204 <= n2572;
/* FF 16 22  1 */ always @(posedge n3) if (n881) io_33_30_1 <= 1'b0 ? 1'b0 : n2573;
/* FF 13 21  0 */ assign io_0_22_0 = n2574;
/* FF 20 18  6 */ always @(posedge n3, posedge n5) if (n5) n1482 <= 1'b0; else if (n1369) n1482 <= n2575;
/* FF 20 15  5 */ assign n1117 = n2576;
/* FF 11 13  7 */ always @(posedge n3, posedge n5) if (n5) n304 <= 1'b0; else if (n441) n304 <= n2577;
/* FF 13  7  1 */ assign n2578 = n655;
/* FF 15 25  0 */ always @(posedge n3, posedge n5) if (n5) n893 <= 1'b0; else if (n2) n893 <= n2579;
/* FF 15 20  7 */ assign n860 = n2580;
/* FF 18 11  3 */ always @(posedge n3, posedge n5) if (n5) n1162 <= 1'b0; else if (n1179) n1162 <= n2581;
/* FF 12 17  6 */ always @(posedge n3) if (1'b1) n490 <= n128 ? 1'b0 : n2582;
/* FF 17 17  2 */ assign n1106 = n2583;
/* FF 22 23  2 */ always @(posedge n3, posedge n5) if (n5) n1700 <= 1'b0; else if (n1656) n1700 <= n2584;
/* FF 11  9  4 */ assign n277 = n2585;
/* FF 16 21  0 */ always @(posedge n3, posedge n5) if (n5) n998 <= 1'b0; else if (n995) n998 <= n2586;
/* FF 13 22  1 */ assign n633 = n2587;
/* FF 20 17  7 */ always @(posedge n3, posedge n5) if (n5) n1474 <= 1'b0; else if (n793) n1474 <= n2588;
/* FF 20 14  6 */ assign n1447 = n2589;
/* FF 23 20  5 */ always @(posedge n3, posedge n5) if (n5) n1508 <= 1'b0; else if (n1655) n1508 <= n2590;
/* FF 14 18  0 */ always @(posedge n3, posedge n5) if (n5) n385 <= 1'b0; else if (1'b1) n385 <= n2591;
/* FF 17 18  3 */ assign n2592 = n2593;
/* FF 21 22  2 */ assign n1564 = n2594;
/* FF 11 22  5 */ always @(posedge n3, posedge n5) if (n5) n403 <= 1'b0; else if (n273) n403 <= n2595;
/* FF 16 15  6 */ assign n802 = n1099;
/* FF 10 15  6 */ always @(posedge n1) if (1'b1) n225 <= n7 ? 1'b0 : n2596;
/* FF 16 20  7 */ assign n996 = n2597;
/* FF 21 24  1 */ always @(posedge n3) if (n688) n1621 <= 1'b0 ? 1'b0 : n2598;
/* FF 15 18  4 */ always @(posedge n3, posedge n5) if (n5) n821 <= 1'b0; else if (n826) n821 <= n2599;
/* FF 18 14  1 */ assign n1190 = n2600;
/* FF 20 16  0 */ always @(posedge n3, posedge n5) if (n5) n1442 <= 1'b0; else if (n1455) n1442 <= n2601;
/* FF 12 20  6 */ always @(posedge n3, posedge n5) if (n5) n522 <= 1'b0; else if (n538) n522 <= n2602;
/* FF 20 13  7 */ always @(posedge n3, posedge n5) if (n5) n1441 <= 1'b0; else if (n933) n1441 <= n2603;
/* FF 11 11  5 */ always @(posedge n1, posedge n5) if (n5) n281 <= 1'b0; else if (1'b1) n281 <= n2604;
/* FF 22 18  2 */ always @(posedge n1, posedge n5) if (n5) n1047 <= 1'b0; else if (n8) n1047 <= n2605;
/* FF  9 15  4 */ assign n162 = n2606;
/* FF 21 10  5 */ assign n1537 = n1630;
/* FF 12 23  0 */ assign n2607 = n2608;
/* FF 14 13  1 */ always @(posedge n3, posedge n5) if (n5) n217 <= 1'b0; else if (n690) n217 <= n2609;
/* FF 19 22  2 */ always @(posedge n3, posedge n5) if (n5) n1391 <= 1'b0; else if (1'b1) n1391 <= n2610;
/* FF 22 17  4 */ assign n2611 = n1732;
/* FF 16 16  4 */ always @(posedge n3, posedge n5) if (n5) n965 <= 1'b0; else if (n799) n965 <= n2612;
/* FF  7 12  2 */ assign n111 = n2613;
/* FF 15 13  2 */ assign n441 = n2614;
/* FF 20 20  5 */ always @(posedge n3, posedge n5) if (n5) n1257 <= 1'b0; else if (n996) n1257 <= n2615;
/* FF 16 14  5 */ assign n948 = n1086;
/* FF 16 19  6 */ always @(posedge n3, posedge n5) if (n5) n991 <= 1'b0; else if (n801) n991 <= n2616;
/* FF 15 19  7 */ always @(posedge n3, posedge n5) if (n5) n842 <= 1'b1; else if (n629) n842 <= n2617;
/* FF 18 17  0 */ assign n1215 = n2618;
/* FF 15 14  4 */ always @(posedge n3, posedge n5) if (n5) n770 <= 1'b0; else if (1'b1) n770 <= n2619;
/* FF 19  9  0 */ always @(posedge n3, posedge n5) if (n5) n1164 <= 1'b0; else if (n596) n1164 <= n2620;
/* FF 21 11  2 */ always @(posedge n3, posedge n5) if (n5) n1542 <= 1'b0; else if (n1631) n1542 <= n2621;
/* FF 18 12  6 */ always @(posedge n3, posedge n5) if (n5) n1175 <= 1'b0; else if (n1298) n1175 <= n2622;
/* FF 12 22  3 */ assign n2623 = n2624;
/* FF 14 12  2 */ assign n676 = n2625;
/* FF 19 23  1 */ always @(posedge n3, posedge n5) if (n5) n1400 <= 1'b0; else if (1'b1) n1400 <= n2626;
/* FF 22 16  7 */ assign n1662 = n2627;
/* FF 20 11  4 */ always @(posedge n3, posedge n5) if (n5) n1430 <= 1'b0; else if (n1199) n1430 <= n2628;
/* FF 19 24  5 */ always @(posedge n3, posedge n5) if (n5) n1410 <= 1'b0; else if (n1025) n1410 <= n2629;
/* FF 11 20  7 */ assign n394 = n2630;
/* FF 16 13  4 */ assign n936 = n2631;
/* FF 16 18  5 */ always @(posedge n3, posedge n5) if (n5) n844 <= 1'b0; else if (n800) n844 <= n2632;
/* FF 15 16  6 */ assign n141 = n972;
/* FF 21 15  7 */ always @(posedge n3, posedge n5) if (n5) n1576 <= 1'b0; else if (n933) n1576 <= n2633;
/* FF 15 15  7 */ always @(posedge n3, posedge n5) if (n5) n791 <= 1'b0; else if (n944) n791 <= n2634;
/* FF 18 16  3 */ always @(posedge n1, posedge n5) if (n5) n705 <= 1'b0; else if (n8) n705 <= n2635;
/* FF 20 22  2 */ always @(posedge n3, posedge n5) if (n5) n1504 <= 1'b0; else if (1'b1) n1504 <= n2636;
/* FF 17 24  0 */ assign n2637 = n2638;
/* FF 24 15  2 */ always @(posedge n3, posedge n5) if (n5) n1602 <= 1'b0; else if (n958) n1602 <= n2639;
/* FF 13 11  5 */ always @(posedge io_0_6_1, posedge n5) if (n5) n562 <= 1'b0; else if (1'b1) n562 <= n2640;
/* FF 21 12  3 */ always @(posedge n3, posedge n5) if (n5) n1548 <= 1'b0; else if (n1186) n1548 <= n2641;
/* FF 12 21  2 */ assign n532 = n2642;
/* FF 19 20  0 */ always @(posedge n3, posedge n5) if (n5) n1376 <= 1'b0; else if (1'b1) n1376 <= n2643;
/* FF 22 19  6 */ assign n1350 = n2644;
/* FF 23 16  4 */ always @(posedge n3, posedge n5) if (n5) n1597 <= 1'b0; else if (n1653) n1597 <= n2645;
/* FF 11 21  0 */ assign n258 = n2646;
/* FF 16 12  3 */ assign n2647 = n1071;
/* FF 16 17  4 */ always @(posedge n3, posedge n5) if (n5) n825 <= 1'b0; else if (n702) n825 <= n2648;
/* FF 13 15  2 */ always @(posedge n3) if (io_0_25_1) n579 <= 1'b0 ? 1'b0 : n2649;
/* FF 15 17  1 */ always @(posedge n3, posedge n5) if (n5) n809 <= 1'b0; else if (n609) n809 <= n2650;
/* FF 18 19  2 */ assign n1230 = n2651;
/* FF 20 21  3 */ always @(posedge n3, posedge n5) if (n5) n1497 <= 1'b0; else if (n1012) n1497 <= n2652;
/* FF 17 25  3 */ assign n1149 = n2653;
/* FF 23 13  1 */ always @(posedge n3, posedge n5) if (n5) n1710 <= 1'b0; else if (n793) n1710 <= n2654;
/* FF 24 14  1 */ always @(posedge n3, posedge n5) if (n5) n1422 <= 1'b0; else if (n467) n1422 <= n2655;
/* FF 13 12  4 */ always @(posedge io_0_6_1, posedge n5) if (n5) n568 <= 1'b0; else if (1'b1) n568 <= n2656;
/* FF 21 13  0 */ assign n1551 = n2657;
/* FF 17 11  0 */ assign n1057 = n2658;
/* FF 19 21  7 */ always @(posedge n3, posedge n5) if (n5) n1286 <= 1'b0; else if (n1145) n1286 <= n2659;
/* FF 11 17  5 */ assign n356 = n2660;
/* FF 23 14  5 */ always @(posedge n3, posedge n5) if (n5) n1718 <= 1'b0; else if (n127) n1718 <= n2661;
/* FF 24 17  5 */ always @(posedge n3, posedge n5) if (n5) n1240 <= 1'b0; else if (n1454) n1240 <= n2662;
/* FF 15 21  6 */ assign n875 = n2663;
/* FF 12 10  2 */ assign n2664 = n556;
/* FF 23 17  3 */ assign n2665 = n1746;
/* FF 11 18  1 */ assign n367 = n2666;
/* FF 16 11  2 */ always @(posedge n3, posedge n5) if (n5) n925 <= 1'b0; else if (n938) n925 <= n2667;
/* FF 13 16  3 */ always @(posedge n3, posedge n5) if (n5) n585 <= 1'b0; else if (n492) n585 <= n2668;
/* FF 15 22  0 */ assign n2669 = n2670;
/* FF 18  9  4 */ always @(posedge n3, posedge n5) if (n5) n917 <= 1'b0; else if (n215) n917 <= n2671;
/* FF 18 18  5 */ assign n2672 = n1364;
/* FF  6 11  3 */ always @(posedge n1, posedge n5) if (n5) n70 <= 1'b0; else if (1'b1) n70 <= n2673;
/* FF 14 10  1 */ always @(posedge n1, posedge n5) if (n5) n659 <= 1'b0; else if (n672) n659 <= n2674;
/* FF 19 17  4 */ assign n2675 = n1478;
/* FF 22 21  7 */ always @(posedge n3, posedge n5) if (n5) n1227 <= 1'b0; else if (n1652) n1227 <= n2676;
/* FF  5 17  2 */ always @(posedge n3, posedge n5) if (n5) n17 <= 1'b0; else if (n4) n17 <= n2677;
/* FF 24 13  0 */ always @(posedge n3, posedge n5) if (n5) n1577 <= 1'b0; else if (n805) n1577 <= n2678;
/* FF 21 14  1 */ assign n1092 = n2679;
/* FF  9 16  2 */ assign n167 = n2680;
/* FF 14 20  6 */ always @(posedge n3, posedge n5) if (n5) n190 <= 1'b0; else if (1'b1) n190 <= n2681;
/* FF 14  9  5 */ assign n411 = n2682;
/* FF 17 20  1 */ assign n1120 = n2683;
/* FF 19 18  6 */ assign n1358 = n2684;
/* FF 10 10  2 */ assign n198 = n2685;
/* FF 23 15  6 */ always @(posedge n3, posedge n5) if (n5) n942 <= 1'b0; else if (n1654) n942 <= n2686;
/* FF 21 16  0 */ always @(posedge n3, posedge n5) if (n5) n1579 <= 1'b0; else if (n596) n1579 <= n2687;
/* FF 15 10  7 */ always @(posedge n1, posedge n5) if (n5) n749 <= 1'b0; else if (1'b1) n749 <= n2688;
/* FF 12  9  3 */ assign n406 = n2689;
/* FF 18 22  2 */ assign n1025 = n1399;
/* FF 11 19  2 */ assign n377 = n2690;
/* FF  9 12  4 */ assign n155 = n2691;
/* FF 13 17  0 */ assign n179 = n2692;
/* FF 18 21  4 */ always @(posedge n3) if (n881) io_33_4_1 <= 1'b0 ? 1'b0 : n2693;
/* FF 19 14  5 */ assign n1311 = n2694;
/* FF 22 20  4 */ assign n1672 = n2695;
/* FF 10 14  7 */ assign n216 = n2696;
/* FF  5 18  3 */ always @(posedge n3, posedge n5) if (n5) n55 <= 1'b0; else if (n4) n55 <= n2697;
/* FF 16 24  5 */ always @(posedge n3, posedge n5) if (n5) n146 <= 1'b0; else if (n1010) n146 <= n2698;
/* FF  9 17  1 */ always @(posedge n3, posedge n5) if (n5) n173 <= 1'b0; else if (n172) n173 <= n2699;
/* FF 14 23  7 */ always @(posedge n3, posedge n5) if (n5) n539 <= 1'b1; else if (n538) n539 <= n2700;
/* FF 20 12  6 */ always @(posedge n3, posedge n5) if (n5) n1103 <= 1'b0; else if (n1299) n1103 <= n2701;
/* FF 19 19  5 */ always @(posedge n3, posedge n5) if (n5) n1078 <= 1'b0; else if (n985) n1078 <= n2702;
/* FF 10 13  3 */ always @(posedge n1, posedge n5) if (n5) n208 <= 1'b0; else if (n138) n208 <= n2703;
/* FF 23 12  7 */ always @(posedge n3) if (n1301) n795 <= 1'b0 ? 1'b0 : n2704;
/* FF 21 17  3 */ always @(posedge n3, posedge n5) if (n5) n1587 <= 1'b0; else if (n1179) n1587 <= n2705;
/* FF 15 11  4 */ always @(posedge n1, posedge n5) if (n5) n763 <= 1'b0; else if (1'b1) n763 <= n2706;
/* FF 18 25  3 */ assign n1276 = n2707;
/* FF 20 15  0 */ assign n1453 = n2708;
/* FF 11 16  3 */ always @(posedge n3, posedge n5) if (n5) n340 <= 1'b0; else if (1'b1) n340 <= n2709;
/* FF 16  9  0 */ always @(posedge n3, posedge n5) if (n5) n913 <= 1'b0; else if (n933) n913 <= n2710;
/* FF 13 18  1 */ assign n182 = n2711;
/* FF 15 20  2 */ assign n855 = n2712;
/* FF 18 20  7 */ assign n1239 = n2713;
/* FF 16  7  3 */ always @(negedge io_0_6_1, posedge n5) if (n5) n903 <= 1'b0; else if (1'b1) n903 <= n2714;
/* FF 19 15  6 */ assign n2715 = n1465;
/* FF 22 23  5 */ always @(posedge n3, posedge n5) if (n5) n1418 <= 1'b0; else if (n1656) n1418 <= n2716;
/* FF 15 26  1 */ always @(posedge n3, posedge n5) if (n5) n899 <= 1'b0; else if (n2) n899 <= n2717;
/* FF  9 18  0 */ always @(posedge n3, posedge n5) if (n5) n176 <= 1'b0; else if (n172) n176 <= n2718;
/* FF 12 12  1 */ always @(posedge io_0_6_1, posedge n5) if (n5) n424 <= 1'b0; else if (n563) n424 <= n2719;
/* FF 14 22  0 */ always @(posedge n3, posedge n5) if (n5) n722 <= 1'b0; else if (n704) n722 <= n2720;
/* FF 17 22  3 */ assign n1132 = n2721;
/* FF 14 11  7 */ always @(posedge n1, posedge n5) if (n5) n671 <= 1'b0; else if (1'b1) n671 <= n2722;
/* FF 19 16  4 */ always @(posedge n3, posedge n5) if (n5) n1337 <= 1'b0; else if (n949) n1337 <= n2723;
/* FF 22 10  0 */ assign n2724 = n2725;
/* FF 21 18  2 */ always @(posedge n3, posedge n5) if (n5) n1593 <= 1'b0; else if (n958) n1593 <= n2727;
/* FF 12 15  5 */ assign n464 = n2728;
/* FF 15  7  4 */ assign n737 = n2729;
/* FF 20 14  3 */ assign n2730 = n1569;
/* FF 23 20  0 */ always @(posedge n3, posedge n5) if (n5) n1228 <= 1'b0; else if (n1655) n1228 <= n2731;
/* FF 13 19  6 */ assign n524 = n2732;
/* FF 18 23  6 */ always @(posedge n3) if (n881) io_33_4_0 <= 1'b0 ? 1'b0 : n2733;
/* FF 14 18  5 */ always @(posedge n3, posedge n5) if (n5) n345 <= 1'b0; else if (1'b1) n345 <= n2734;
/* FF 14  7  2 */ always @(negedge io_0_6_1, posedge n5) if (n5) n648 <= 1'b0; else if (1'b1) n648 <= n2735;
/* FF 19 12  7 */ assign n157 = n2736;
/* FF 12 19  0 */ always @(posedge n3, posedge n5) if (n5) n503 <= 1'b0; else if (n620) n503 <= n2737;
/* FF 14 17  1 */ assign n707 = n2738;
/* FF 17 12  5 */ assign n1067 = n2739;
/* FF 17 23  4 */ assign n1141 = n2740;
/* FF 10 15  1 */ always @(posedge n1) if (1'b1) n220 <= n7 ? 1'b0 : n2741;
/* FF 21 19  5 */ assign n2742 = n1684;
/* FF 13 23  3 */ assign n2743 = n2744;
/* FF 18 14  6 */ always @(posedge n1, posedge n5) if (n5) n1053 <= 1'b0; else if (n8) n1053 <= n2745;
/* FF 15  9  2 */ always @(posedge n3, posedge n5) if (n5) n746 <= 1'b0; else if (1'b1) n746 <= n2746;
/* FF 12 14  6 */ assign n448 = n2747;
/* FF 20 13  2 */ assign n1437 = n2748;
/* FF 10 17  5 */ always @(posedge n1) if (1'b1) n228 <= n7 ? 1'b0 : n2749;
/* FF  9 15  1 */ assign n161 = n2750;
/* FF 13 20  7 */ assign n628 = n2751;
/* FF 18 13  0 */ assign n2752 = n1312;
/* FF 20 19  1 */ always @(posedge n3, posedge n5) if (n5) n1490 <= 1'b0; else if (n803) n1490 <= n2753;
/* FF 14 13  4 */ always @(posedge n3, posedge n5) if (n5) n686 <= 1'b0; else if (n690) n686 <= n2754;
/* FF 17 19  1 */ assign n2755 = n2756;
/* FF 19 13  0 */ always @(posedge n3, posedge n5) if (n5) n1303 <= 1'b0; else if (n596) n1303 <= n2757;
/* FF 22 17  3 */ assign n1667 = n2758;
/* FF 15 24  3 */ always @(posedge n3, posedge n5) if (n5) n887 <= 1'b0; else if (n2) n887 <= n2759;
/* FF 21 23  2 */ always @(posedge n3, posedge n5) if (n5) n1282 <= 1'b0; else if (n1453) n1282 <= n2760;
/* FF 15 13  7 */ always @(posedge n3, posedge n5) if (n5) n779 <= 1'b0; else if (n321) n779 <= n2761;
/* FF 12 18  3 */ always @(posedge n3) if (1'b1) n487 <= n128 ? 1'b0 : n2762;
/* FF 14 16  2 */ always @(posedge n3, posedge n5) if (n5) n699 <= 1'b0; else if (1'b1) n699 <= n2763;
/* FF 17 13  6 */ assign n2764 = n1189;
/* FF 17 16  5 */ assign n2765 = n1214;
/* FF 21 20  4 */ always @(posedge n3, posedge n5) if (n5) n1605 <= 1'b0; else if (n270) n1605 <= n2766;
/* FF 13 24  2 */ assign n2767 = n2768;
/* FF 15 14  3 */ assign n540 = n2769;
/* FF 18 17  7 */ assign n1218 = n2770;
/* FF 12 13  7 */ always @(posedge n3, posedge n5) if (n5) n438 <= 1'b0; else if (n573) n438 <= n2771;
/* FF 10 16  6 */ always @(posedge n1) if (1'b1) n236 <= n7 ? 1'b0 : n2772;
/* FF 18 12  3 */ always @(posedge n3, posedge n5) if (n5) n1172 <= 1'b0; else if (n1298) n1172 <= n2773;
/* FF 20 18  2 */ assign n934 = n2774;
/* FF 19 10  1 */ always @(posedge n3, posedge n5) if (n5) n1163 <= 1'b0; else if (n580) n1163 <= n2775;
/* FF 22 16  0 */ always @(posedge n3, posedge n5) if (n5) n1659 <= 1'b0; else if (n596) n1659 <= n2776;
/* FF 15 25  4 */ always @(posedge n3, posedge n5) if (n5) n541 <= 1'b0; else if (n2) n541 <= n2777;
/* FF 12 17  2 */ always @(posedge n3) if (1'b1) n470 <= n128 ? 1'b0 : n2778;
/* FF 14 19  3 */ always @(posedge n3, posedge n5) if (n5) n514 <= 1'b0; else if (1'b1) n514 <= n2779;
/* FF 17 14  7 */ assign n1083 = n2780;
/* FF 19 24  0 */ always @(posedge n3, posedge n5) if (n5) n1405 <= 1'b0; else if (n1025) n1405 <= n2781;
/* FF 17 17  6 */ assign n1109 = n2782;
/* FF 21 21  7 */ assign n1614 = n2783;
/* FF 15 15  0 */ always @(posedge n3, posedge n5) if (n5) n483 <= 1'b0; else if (n944) n483 <= n2784;
/* FF 18 16  4 */ always @(posedge n1, posedge n5) if (n5) n1180 <= 1'b0; else if (n8) n1180 <= n2785;
/* FF 10 19  7 */ always @(posedge n3, posedge n5) if (n5) n254 <= 1'b0; else if (n359) n254 <= n2786;
/* FF 13 11  2 */ always @(posedge io_0_6_1, posedge n5) if (n5) n559 <= 1'b0; else if (1'b1) n559 <= n2787;
/* FF 13 22  5 */ assign n637 = n2788;
/* FF 18 15  2 */ assign n2789 = n1333;
/* FF  6 12  2 */ assign n77 = n2790;
/* FF 20 17  3 */ always @(posedge n3, posedge n5) if (n5) n1470 <= 1'b0; else if (n793) n1470 <= n2791;
/* FF 14 15  6 */ assign n321 = n2792;
/* FF 19 11  2 */ always @(posedge n3, posedge n5) if (n5) n1296 <= 1'b0; else if (n1300) n1296 <= n2793;
/* FF 22 19  1 */ always @(posedge n3, posedge n5) if (n5) n1615 <= 1'b0; else if (n1369) n1615 <= n2794;
/* FF 12 16  5 */ assign n482 = n2795;
/* FF 17 15  0 */ assign n2796 = n1205;
/* FF 17 18  7 */ assign n2797 = n2798;
/* FF 22 13  5 */ always @(posedge n3, posedge n5) if (n5) n1641 <= 1'b0; else if (n805) n1641 <= n2799;
/* FF 15 12  1 */ always @(posedge n3, posedge n5) if (n5) n358 <= 1'b0; else if (1'b1) n358 <= n2800;
/* FF 18 19  5 */ assign n1236 = n2801;
/* FF 11 22  1 */ always @(posedge n3, posedge n5) if (n5) n399 <= 1'b0; else if (n273) n399 <= n2802;
/* FF 16 15  2 */ assign n702 = n2803;
/* FF 10 18  0 */ always @(posedge n1) if (n153) n239 <= n7 ? 1'b0 : n2804;
/* FF 13 12  3 */ always @(posedge io_0_6_1, posedge n5) if (n5) n567 <= 1'b0; else if (1'b1) n567 <= n2805;
/* FF 15 18  0 */ always @(posedge n3, posedge n5) if (n5) n815 <= 1'b0; else if (n826) n815 <= n2806;
/* FF 20 16  4 */ always @(posedge n3, posedge n5) if (n5) n1468 <= 1'b0; else if (n1455) n1468 <= n2807;
/* FF 12 20  2 */ always @(posedge n3, posedge n5) if (n5) n519 <= 1'b0; else if (n538) n519 <= n2808;
/* FF 14 14  1 */ assign n32 = n2809;
/* FF 17 11  5 */ assign n1060 = n2810;
/* FF 19  8  3 */ always @(posedge n1, posedge n5) if (n5) n931 <= 1'b0; else if (n672) n931 <= n2811;
/* FF 23 14  0 */ always @(posedge n3, posedge n5) if (n5) n1461 <= 1'b0; else if (n127) n1461 <= n2812;
/* FF 24 17  0 */ always @(posedge n3, posedge n5) if (n5) n1591 <= 1'b0; else if (n1454) n1591 <= n2813;
/* FF 21 10  1 */ assign n8 = n2814;
/* FF 12 10  7 */ assign n410 = n2815;
/* FF 12 23  4 */ assign n2816 = n2817;
/* FF 17  8  1 */ always @(posedge n3, posedge n5) if (n5) n910 <= 1'b0; else if (1'b1) n910 <= n2818;
/* FF 16 16  0 */ always @(posedge n3, posedge n5) if (n5) n814 <= 1'b0; else if (n799) n814 <= n2819;
/* FF 22 12  6 */ always @(posedge n3, posedge n5) if (n5) n804 <= 1'b0; else if (n1077) n804 <= n2820;
/* FF 13 16  6 */ always @(posedge n3, posedge n5) if (n5) n588 <= 1'b0; else if (n492) n588 <= n2821;
/* FF  7 12  6 */ assign n121 = n137;
/* FF 18 18  2 */ assign n1223 = n2822;
/* FF 20 20  1 */ always @(posedge n3, posedge n5) if (n5) n1493 <= 1'b0; else if (n996) n1493 <= n2823;
/* FF 23 18  2 */ always @(posedge n3, posedge n5) if (n5) n1734 <= 1'b0; else if (n1117) n1734 <= n2824;
/* FF 16 14  1 */ assign n467 = n2825;
/* FF  5 17  7 */ always @(posedge n3, posedge n5) if (n5) n27 <= 1'b0; else if (n4) n27 <= n2826;
/* FF 13 13  0 */ always @(posedge io_0_6_1, posedge n5) if (n5) n571 <= 1'b0; else if (n563) n571 <= n2827;
/* FF 15 19  3 */ always @(posedge n3, posedge n5) if (n5) n838 <= 1'b1; else if (n629) n838 <= n2828;
/* FF 20 23  5 */ always @(posedge n3) if (n688) n1520 <= 1'b0 ? 1'b0 : n2829;
/* FF 14  9  0 */ assign n657 = n2830;
/* FF 17 20  4 */ assign n1123 = n2831;
/* FF 23 15  3 */ always @(posedge n3, posedge n5) if (n5) n1719 <= 1'b0; else if (n1654) n1719 <= n2832;
/* FF 21 16  7 */ assign n1582 = n2833;
/* FF 21 11  6 */ always @(posedge n3, posedge n5) if (n5) n430 <= 1'b0; else if (n1631) n430 <= n2834;
/* FF 18 22  7 */ always @(posedge n3, posedge n5) if (n5) n1021 <= 1'b0; else if (1'b1) n1021 <= n2835;
/* FF 12 22  7 */ assign n2836 = n2837;
/* FF 10  9  3 */ always @(posedge n1, posedge n5) if (n5) n196 <= 1'b0; else if (1'b1) n196 <= n2838;
/* FF 22 15  7 */ assign n1656 = n2839;
/* FF 13 17  5 */ assign n246 = n2840;
/* FF 18 21  3 */ always @(posedge n3) if (n881) io_20_33_1 <= 1'b0 ? 1'b0 : n2841;
/* FF 20 11  0 */ always @(posedge n3, posedge n5) if (n5) n1427 <= 1'b0; else if (n1199) n1427 <= n2842;
/* FF 23 19  1 */ assign n1735 = n2843;
/* FF 11 20  3 */ assign n390 = n2844;
/* FF 16 13  0 */ assign n690 = n2845;
/* FF  5 18  6 */ always @(posedge n3, posedge n5) if (n5) n58 <= 1'b0; else if (n4) n58 <= n2846;
/* FF 10 20  2 */ always @(posedge n3, posedge n5) if (n5) n261 <= 1'b0; else if (n144) n261 <= n2847;
/* FF 15 16  2 */ assign n799 = n2848;
/* FF 21 15  3 */ assign n2849 = n1658;
/* FF 20 25  7 */ always @(posedge n3, posedge n5) if (n5) n1420 <= 1'b0; else if (n1453) n1420 <= n2850;
/* FF 20 22  6 */ always @(posedge n3, posedge n5) if (n5) io_11_33_1 <= 1'b0; else if (1'b1) io_11_33_1 <= n2851;
/* FF 17 24  4 */ assign n2852 = n2853;
/* FF 23 12  2 */ always @(posedge n3) if (n1301) n1608 <= 1'b0 ? 1'b0 : n2854;
/* FF  7 10  7 */ always @(posedge n1, posedge n5) if (n5) io_4_0_0 <= 1'b0; else if (1'b1) io_4_0_0 <= n2855;
/* FF 21 17  4 */ assign n1475 = n2856;
/* FF 21 12  7 */ always @(posedge n3, posedge n5) if (n5) n1194 <= 1'b0; else if (n1186) n1194 <= n2857;
/* FF 18 25  6 */ assign n1279 = n2858;
/* FF 12 21  6 */ assign n536 = n2859;
/* FF 22 14  0 */ always @(posedge n3, posedge n5) if (n5) n1434 <= 1'b0; else if (n1651) n1434 <= n2860;
/* FF 13 18  4 */ assign n605 = n2861;
/* FF 18 20  0 */ assign n2862 = n1385;
/* FF 20 10  3 */ always @(posedge n1, posedge n5) if (n5) n1425 <= 1'b0; else if (1'b1) n1425 <= n2863;
/* FF 23 16  0 */ always @(posedge n3, posedge n5) if (n5) n439 <= 1'b0; else if (n1653) n439 <= n2864;
/* FF 11 14  5 */ assign n317 = n2865;
/* FF 16 12  7 */ assign n703 = n2866;
/* FF  5 19  1 */ always @(posedge n3, posedge n5) if (n5) n61 <= 1'b0; else if (n4) n61 <= n2867;
/* FF 22 24  1 */ always @(posedge n3, posedge n5) if (n5) n1417 <= 1'b0; else if (n1369) n1417 <= n2868;
/* FF 15 17  5 */ always @(posedge n3, posedge n5) if (n5) n714 <= 1'b0; else if (n609) n714 <= n2869;
/* FF 12 12  6 */ always @(posedge io_0_6_1, posedge n5) if (n5) n428 <= 1'b0; else if (n563) n428 <= n2870;
/* FF 20 21  7 */ always @(posedge n3, posedge n5) if (n5) n1499 <= 1'b0; else if (n1012) n1499 <= n2871;
/* FF 17 22  6 */ assign n1135 = n2872;
/* FF 14 11  2 */ always @(posedge n1, posedge n5) if (n5) n667 <= 1'b0; else if (1'b1) n667 <= n2873;
/* FF 22 10  5 */ assign n1625 = n2874;
/* FF 21 18  5 */ always @(posedge n3, posedge n5) if (n5) n1595 <= 1'b0; else if (n958) n1595 <= n2875;
/* FF 21 13  4 */ always @(posedge n3, posedge n5) if (n5) n1553 <= 1'b0; else if (n596) n1553 <= n2876;
/* FF 12 15  0 */ assign n459 = n2877;
/* FF 15  7  1 */ assign n734 = n906;
/* FF 18 24  5 */ assign n816 = n2878;
/* FF 11 17  1 */ assign n128 = n2879;
/* FF 13 19  3 */ assign n131 = n2880;
/* FF 15 21  2 */ assign n871 = n2881;
/* FF 18 23  1 */ always @(posedge n3) if (n881) io_33_29_1 <= 1'b0 ? 1'b0 : n2882;
/* FF 23 17  7 */ assign n608 = n2883;
/* FF 11 15  6 */ assign n329 = n2884;
/* FF 14  7  5 */ always @(negedge io_0_6_1, posedge n5) if (n5) n651 <= 1'b0; else if (1'b1) n651 <= n2885;
/* FF 11 18  5 */ assign n371 = n2886;
/* FF 16 11  6 */ always @(posedge n3, posedge n5) if (n5) n927 <= 1'b0; else if (n938) n927 <= n2887;
/* FF 15 22  4 */ assign n2888 = n2889;
/* FF 18  9  0 */ always @(posedge n3, posedge n5) if (n5) n1155 <= 1'b0; else if (n215) n1155 <= n2890;
/* FF 12 19  7 */ always @(posedge n3, posedge n5) if (n5) n510 <= 1'b1; else if (n620) n510 <= n2891;
/* FF  6 11  7 */ always @(posedge n1, posedge n5) if (n5) n74 <= 1'b0; else if (1'b1) n74 <= n2892;
/* FF 17 23  1 */ assign n1138 = n2893;
/* FF 19 17  0 */ assign n2894 = n1476;
/* FF 22 21  3 */ always @(posedge n3, posedge n5) if (n5) n1693 <= 1'b0; else if (n1652) n1693 <= n2895;
/* FF  7  8  5 */ always @(posedge n1, posedge n5) if (n5) io_4_0_1 <= 1'b1; else if (1'b1) io_4_0_1 <= n2896;
/* FF 21 19  2 */ assign n1601 = n2897;
/* FF 21 14  5 */ always @(posedge n3, posedge n5) if (n5) n1561 <= 1'b0; else if (n805) n1561 <= n2898;
/* FF 12 14  3 */ assign n445 = n2899;
/* FF 14 20  2 */ always @(posedge n3, posedge n5) if (n5) n528 <= 1'b0; else if (1'b1) n528 <= n2900;
/* FF 10 10  6 */ assign n2901 = n2902;
/* FF 16 23  5 */ always @(posedge n3, posedge n5) if (n5) n1019 <= 1'b0; else if (n1010) n1019 <= n2903;
/* FF 13 20  2 */ assign n623 = n2904;
/* FF 20 19  4 */ always @(posedge n3, posedge n5) if (n5) n1256 <= 1'b0; else if (n803) n1256 <= n2905;
/* FF 11 12  7 */ always @(posedge n3, posedge n5) if (n5) n218 <= 1'b0; else if (n26) n218 <= n2906;
/* FF 17 19  6 */ assign n2907 = n2908;
/* FF 11 19  6 */ assign n381 = n2909;
/* FF 16 10  5 */ always @(posedge n1, posedge n5) if (n5) n669 <= 1'b0; else if (n672) n669 <= n2910;
/* FF 15 24  6 */ always @(posedge n3, posedge n5) if (n5) n890 <= 1'b0; else if (n2) n890 <= n2911;
/* FF 12 18  4 */ always @(posedge n3) if (1'b1) n499 <= n128 ? 1'b0 : n2912;
/* FF 17 16  0 */ assign n1100 = n2913;
/* FF 19 14  1 */ assign n2914 = n1450;
/* FF 22 20  0 */ assign n1679 = n2915;
/* FF 10 14  3 */ assign n215 = n2916;
/* FF 16 24  1 */ always @(posedge n3, posedge n5) if (n5) n543 <= 1'b0; else if (n1010) n543 <= n2917;
/* FF 21 20  3 */ always @(posedge n3, posedge n5) if (n5) n1604 <= 1'b0; else if (n270) n1604 <= n2918;
/* FF  9 17  5 */ always @(posedge n3, posedge n5) if (n5) n174 <= 1'b0; else if (n172) n174 <= n2919;
/* FF 12 13  2 */ always @(posedge n3, posedge n5) if (n5) n433 <= 1'b0; else if (n573) n433 <= n2920;
/* FF 20 12  2 */ always @(posedge n3, posedge n5) if (n5) n1185 <= 1'b0; else if (n1299) n1185 <= n2921;
/* FF 10 13  7 */ always @(posedge n1, posedge n5) if (n5) n211 <= 1'b0; else if (n138) n211 <= n2922;
/* FF 15 11  0 */ always @(posedge n1, posedge n5) if (n5) n761 <= 1'b0; else if (1'b1) n761 <= n2923;
/* FF 20 15  4 */ assign n592 = n1578;
/* FF 11 13  0 */ always @(posedge n3, posedge n5) if (n5) n297 <= 1'b0; else if (n441) n297 <= n2924;
/* FF 11 16  7 */ assign n344 = n2925;
/* FF 13  7  2 */ assign n2926 = n656;
/* FF 15 25  1 */ always @(posedge n3, posedge n5) if (n5) n892 <= 1'b0; else if (n2) n892 <= n2927;
/* FF 18 11  2 */ always @(posedge n3, posedge n5) if (n5) n1161 <= 1'b0; else if (n1179) n1161 <= n2928;
/* FF 15 20  6 */ assign n859 = n2929;
/* FF 12 17  5 */ always @(posedge n3) if (1'b1) n473 <= n128 ? 1'b0 : n2930;
/* FF 17 17  3 */ assign n1107 = n2931;
/* FF 19 15  2 */ assign n1323 = n2932;
/* FF 22 23  1 */ always @(posedge n3, posedge n5) if (n5) n1416 <= 1'b0; else if (n1656) n1416 <= n2933;
/* FF 21 21  0 */ assign n2934 = n1695;
/* FF 14 22  4 */ always @(posedge n3, posedge n5) if (n5) n718 <= 1'b0; else if (n704) n718 <= n2935;
/* FF 11  9  5 */ always @(posedge n1, posedge n5) if (n5) n278 <= 1'b0; else if (1'b1) n278 <= n2936;
/* FF 16 21  7 */ always @(posedge n3, posedge n5) if (n5) n1005 <= 1'b1; else if (n995) n1005 <= n2937;
/* FF 13 22  0 */ assign n632 = n2938;
/* FF 15  8  1 */ assign n544 = n2940;
/* FF 20 17  6 */ assign n1473 = n2941;
/* FF 23 20  4 */ always @(posedge n3, posedge n5) if (n5) n1507 <= 1'b0; else if (n1655) n1507 <= n2942;
/* FF 11 10  1 */ always @(posedge n1, posedge n5) if (n5) n283 <= 1'b0; else if (1'b1) n283 <= n2943;
/* FF  9 14  2 */ always @(posedge n1) if (1'b1) n84 <= 1'b0 ? 1'b0 : n2944;
/* FF 14 18  1 */ always @(posedge n3, posedge n5) if (n5) n256 <= 1'b0; else if (1'b1) n256 <= n2945;
/* FF 17 18  2 */ assign n2946 = n2947;
/* FF 19 12  3 */ assign n1300 = n2948;
/* FF 21 22  1 */ assign n1609 = n2949;
/* FF 14 17  5 */ always @(posedge n1, posedge n5) if (n5) n673 <= 1'b0; else if (n8) n673 <= n2950;
/* FF 17 12  1 */ assign n2951 = n1182;
/* FF 11 22  4 */ always @(posedge n3, posedge n5) if (n5) n402 <= 1'b1; else if (n273) n402 <= n2952;
/* FF 10 15  5 */ always @(posedge n1) if (1'b1) n224 <= n7 ? 1'b0 : n2953;
/* FF 16 20  0 */ always @(posedge n3) if (1'b1) n994 <= 1'b0 ? 1'b0 : n2954;
/* FF 21 24  0 */ always @(posedge n3) if (n688) n1620 <= 1'b0 ? 1'b0 : n2955;
/* FF 15 18  7 */ always @(posedge n3, posedge n5) if (n5) n824 <= 1'b0; else if (n826) n824 <= n2956;
/* FF 18 14  2 */ assign n2957 = n1325;
/* FF 20 16  1 */ always @(posedge n3, posedge n5) if (n5) n1458 <= 1'b0; else if (n1455) n1458 <= n2958;
/* FF 12 20  7 */ always @(posedge n3, posedge n5) if (n5) n523 <= 1'b0; else if (n538) n523 <= n2959;
/* FF 20 13  6 */ assign n1440 = n2960;
/* FF 11 11  2 */ always @(posedge n1, posedge n5) if (n5) n294 <= 1'b0; else if (1'b1) n294 <= n2961;
/* FF 22 18  3 */ assign n1670 = n2962;
/* FF 10 17  1 */ always @(posedge n1) if (1'b1) n240 <= n7 ? 1'b0 : n2963;
/* FF  9 15  5 */ assign n2964 = n230;
/* FF 13  9  0 */ always @(posedge n3, posedge n5) if (n5) n546 <= 1'b0; else if (1'b1) n546 <= n2965;
/* FF 21 10  4 */ assign n2966 = n1629;
/* FF 18 13  4 */ assign n1183 = n2967;
/* FF 12 23  3 */ assign n2968 = n2969;
/* FF 14 13  0 */ always @(posedge n3, posedge n5) if (n5) n683 <= 1'b0; else if (n690) n683 <= n2970;
/* FF 19 22  5 */ always @(posedge n3, posedge n5) if (n5) n1394 <= 1'b0; else if (1'b1) n1394 <= n2971;
/* FF 19 13  4 */ assign n1305 = n2972;
/* FF 16 16  5 */ always @(posedge n3, posedge n5) if (n5) n966 <= 1'b0; else if (n799) n966 <= n2973;
/* FF  7 12  1 */ assign n26 = n2974;
/* FF 15 13  3 */ assign n573 = n2975;
/* FF 20 20  6 */ always @(posedge n3, posedge n5) if (n5) n1118 <= 1'b0; else if (n996) n1118 <= n2976;
/* FF 14 16  6 */ always @(posedge n3, posedge n5) if (n5) n696 <= 1'b0; else if (1'b1) n696 <= n2977;
/* FF 17 13  2 */ assign n1074 = n2978;
/* FF 16 19  1 */ always @(posedge n3, posedge n5) if (n5) n987 <= 1'b0; else if (n801) n987 <= n2979;
/* FF 15 19  4 */ always @(posedge n3, posedge n5) if (n5) n839 <= 1'b1; else if (n629) n839 <= n2980;
/* FF 18 17  3 */ always @(posedge n3, posedge n5) if (n5) n1216 <= 1'b0; else if (n1117) n1216 <= n2981;
/* FF 15 14  7 */ assign n780 = n2982;
/* FF 20 23  0 */ assign n1501 = n2983;
/* FF 10 16  2 */ always @(posedge n1) if (1'b1) n232 <= n7 ? 1'b0 : n2984;
/* FF 13 10  1 */ always @(posedge n1, posedge n5) if (n5) n549 <= 1'b0; else if (1'b1) n549 <= n2985;
/* FF 21 11  3 */ always @(posedge n3, posedge n5) if (n5) n1543 <= 1'b0; else if (n1631) n1543 <= n2986;
/* FF 18 12  7 */ always @(posedge n3, posedge n5) if (n5) n1176 <= 1'b0; else if (n1298) n1176 <= n2987;
/* FF 12 22  0 */ assign n2988 = n2989;
/* FF 14 12  3 */ assign n666 = n2990;
/* FF 19 23  6 */ always @(posedge n3, posedge n5) if (n5) n1404 <= 1'b0; else if (1'b1) n1404 <= n2991;
/* FF 19 10  5 */ always @(posedge n3, posedge n5) if (n5) n1292 <= 1'b0; else if (n580) n1292 <= n2992;
/* FF 22 16  4 */ assign n1661 = n2993;
/* FF 14 19  7 */ always @(posedge n3, posedge n5) if (n5) n513 <= 1'b0; else if (1'b1) n513 <= n2994;
/* FF 17 14  3 */ assign n2995 = n1197;
/* FF 19 24  4 */ always @(posedge n3, posedge n5) if (n5) n1409 <= 1'b0; else if (n1025) n1409 <= n2996;
/* FF 11 20  6 */ assign n393 = n2997;
/* FF 16 18  2 */ always @(posedge n3, posedge n5) if (n5) n980 <= 1'b0; else if (n800) n980 <= n2998;
/* FF 15 16  5 */ assign n800 = n2999;
/* FF 15 15  4 */ always @(posedge n3, posedge n5) if (n5) n788 <= 1'b0; else if (n944) n788 <= n3000;
/* FF 18 16  0 */ assign n3001 = n3002;
/* FF 20 22  3 */ assign n3004 = n1619;
/* FF 17 24  3 */ assign n3005 = n3006;
/* FF 10 19  3 */ always @(posedge n3, posedge n5) if (n5) n250 <= 1'b0; else if (n359) n250 <= n3007;
/* FF 13 11  6 */ assign n563 = n3008;
/* FF 21 12  2 */ always @(posedge n3, posedge n5) if (n5) n1547 <= 1'b0; else if (n1186) n1547 <= n3009;
/* FF 18 15  6 */ assign n1202 = n3010;
/* FF 12 21  1 */ assign n531 = n3011;
/* FF 19 20  7 */ assign n985 = n3012;
/* FF 19 11  6 */ always @(posedge n3, posedge n5) if (n5) n1166 <= 1'b0; else if (n1300) n1166 <= n3013;
/* FF 22 19  5 */ always @(posedge n3, posedge n5) if (n5) n1677 <= 1'b0; else if (n1369) n1677 <= n3014;
/* FF 17 15  4 */ assign n1089 = n3015;
/* FF 16 17  3 */ always @(posedge n3, posedge n5) if (n5) n245 <= 1'b0; else if (n702) n245 <= n3016;
/* FF 22 13  1 */ assign n1638 = n3017;
/* FF 15 17  2 */ always @(posedge n3, posedge n5) if (n5) n810 <= 1'b0; else if (n609) n810 <= n3018;
/* FF 15 12  5 */ always @(posedge n3, posedge n5) if (n5) n125 <= 1'b0; else if (1'b1) n125 <= n3019;
/* FF 18 19  1 */ always @(posedge n3, posedge n5) if (n5) n1233 <= 1'b0; else if (n1117) n1233 <= n3020;
/* FF 20 21  2 */ assign n1495 = n3021;
/* FF 17 25  0 */ assign n712 = n3022;
/* FF 24 14  6 */ always @(posedge n3, posedge n5) if (n5) n792 <= 1'b0; else if (n467) n792 <= n3023;
/* FF 21 13  1 */ assign n3024 = n1643;
/* FF 17 11  1 */ assign n3025 = n1168;
/* FF 19 21  0 */ always @(posedge n3, posedge n5) if (n5) n135 <= 1'b0; else if (n1145) n135 <= n3026;
/* FF 11 17  6 */ assign n3027 = n498;
/* FF 23 14  4 */ always @(posedge n3, posedge n5) if (n5) n1717 <= 1'b0; else if (n127) n1717 <= n3028;
/* FF 24 17  4 */ always @(posedge n3, posedge n5) if (n5) n1744 <= 1'b0; else if (n1454) n1744 <= n3029;
/* FF 15 21  7 */ assign n876 = n3030;
/* FF 12 10  3 */ assign n409 = n3031;
/* FF 17  8  5 */ always @(posedge n3, posedge n5) if (n5) n149 <= 1'b0; else if (1'b1) n149 <= n3032;
/* FF 11 18  0 */ assign n366 = n3033;
/* FF 22 12  2 */ always @(posedge n3, posedge n5) if (n5) n1634 <= 1'b0; else if (n1077) n1634 <= n3035;
/* FF 13 16  2 */ always @(posedge n3, posedge n5) if (n5) n584 <= 1'b0; else if (n492) n584 <= n3036;
/* FF 15 22  3 */ assign n3037 = n3038;
/* FF 18  9  7 */ always @(posedge n3, posedge n5) if (n5) n916 <= 1'b0; else if (n215) n916 <= n3039;
/* FF 18 18  6 */ assign n3040 = n1365;
/* FF  6 11  2 */ always @(posedge n1, posedge n5) if (n5) n69 <= 1'b0; else if (1'b1) n69 <= n3041;
/* FF 14 10  2 */ always @(posedge n1, posedge n5) if (n5) n660 <= 1'b0; else if (n672) n660 <= n3042;
/* FF 19 17  5 */ assign n3043 = n1479;
/* FF 22 21  6 */ always @(posedge n3, posedge n5) if (n5) n1372 <= 1'b0; else if (n1652) n1372 <= n3044;
/* FF  5 17  3 */ always @(posedge n3, posedge n5) if (n5) n47 <= 1'b0; else if (n4) n47 <= n3045;
/* FF 21 14  0 */ assign n3046 = n1648;
/* FF 20 26  2 */ always @(posedge n3, posedge n5) if (n5) n1151 <= 1'b0; else if (n1453) n1151 <= n3047;
/* FF 14 20  7 */ always @(posedge n3, posedge n5) if (n5) n526 <= 1'b0; else if (1'b1) n526 <= n3048;
/* FF 14  9  4 */ assign n3049 = n751;
/* FF 17 20  0 */ assign n1119 = n3050;
/* FF 19 18  1 */ assign n3051 = n1487;
/* FF 10 10  3 */ assign n199 = n3052;
/* FF 23 15  7 */ always @(posedge n3, posedge n5) if (n5) n977 <= 1'b0; else if (n1654) n977 <= n3053;
/* FF 21 16  3 */ assign n3054 = n1664;
/* FF 15 10  6 */ always @(posedge n1, posedge n5) if (n5) n754 <= 1'b0; else if (1'b1) n754 <= n3055;
/* FF 18 22  3 */ assign n1258 = n3056;
/* FF 11 19  3 */ assign n378 = n3057;
/* FF  9 12  7 */ always @(posedge n1, posedge n5) if (n5) n75 <= 1'b0; else if (1'b1) n75 <= n3058;
/* FF 22 15  3 */ assign n1653 = n3059;
/* FF 13 17  1 */ assign n593 = n3060;
/* FF 15 23  0 */ assign n731 = n3061;
/* FF 18 21  7 */ always @(posedge n3) if (n881) io_20_33_0 <= 1'b0 ? 1'b0 : n3062;
/* FF 19 14  4 */ assign n3063 = n1452;
/* FF 22 20  5 */ always @(posedge n3, posedge n5) if (n5) n1686 <= 1'b0; else if (n1117) n1686 <= n3064;
/* FF  5 18  2 */ always @(posedge n3, posedge n5) if (n5) n54 <= 1'b0; else if (n4) n54 <= n3065;
/* FF 16 24  6 */ always @(posedge n3, posedge n5) if (n5) n132 <= 1'b0; else if (n1010) n132 <= n3066;
/* FF 10 20  6 */ always @(posedge n3, posedge n5) if (n5) n265 <= 1'b0; else if (n144) n265 <= n3067;
/* FF 20 25  3 */ always @(posedge n3, posedge n5) if (n5) n1509 <= 1'b0; else if (n1453) n1509 <= n3068;
/* FF 20 12  7 */ always @(posedge n3, posedge n5) if (n5) n1193 <= 1'b0; else if (n1299) n1193 <= n3069;
/* FF 19 19  2 */ always @(posedge n3, posedge n5) if (n5) n1367 <= 1'b0; else if (n985) n1367 <= n3070;
/* FF 10 13  2 */ always @(posedge n1, posedge n5) if (n5) n207 <= 1'b0; else if (n138) n207 <= n3071;
/* FF 23 12  6 */ always @(posedge n3) if (n1301) n953 <= 1'b0 ? 1'b0 : n3072;
/* FF  7 10  3 */ always @(posedge n1, posedge n5) if (n5) n108 <= 1'b1; else if (1'b1) n108 <= n3073;
/* FF 21 17  0 */ assign n1584 = n3074;
/* FF 15 11  5 */ always @(posedge n1, posedge n5) if (n5) n764 <= 1'b0; else if (1'b1) n764 <= n3075;
/* FF 18 25  2 */ assign n1275 = n3076;
/* FF 17  7  0 */ always @(posedge n1, posedge n5) if (n5) n914 <= 1'b0; else if (n8) n914 <= n3077;
/* FF 20 15  3 */ assign n1179 = n3078;
/* FF 17 10  7 */ always @(posedge n1, posedge n5) if (n5) n759 <= 1'b0; else if (n8) n759 <= n3079;
/* FF 22 14  4 */ always @(posedge n3, posedge n5) if (n5) n1341 <= 1'b0; else if (n1651) n1341 <= n3080;
/* FF 13 18  0 */ assign n255 = n3081;
/* FF 15 20  1 */ assign n854 = n3083;
/* FF 18 20  4 */ assign n1246 = n3084;
/* FF 11 14  1 */ assign n313 = n3085;
/* FF 16  7  2 */ always @(negedge io_0_6_1, posedge n5) if (n5) n902 <= 1'b0; else if (1'b1) n902 <= n3086;
/* FF 19 15  7 */ assign n1330 = n3087;
/* FF 22 23  4 */ always @(posedge n3, posedge n5) if (n5) n1421 <= 1'b0; else if (n1656) n1421 <= n3088;
/* FF 15 26  0 */ always @(posedge n3, posedge n5) if (n5) n898 <= 1'b0; else if (n2) n898 <= n3089;
/* FF 12 12  2 */ always @(posedge io_0_6_1, posedge n5) if (n5) n425 <= 1'b0; else if (n563) n425 <= n3090;
/* FF 17 22  2 */ assign n1131 = n3091;
/* FF 14 11  6 */ always @(posedge n1, posedge n5) if (n5) n665 <= 1'b0; else if (1'b1) n665 <= n3092;
/* FF 19 16  3 */ always @(posedge n3, posedge n5) if (n5) n1336 <= 1'b0; else if (n949) n1336 <= n3093;
/* FF 10 12  1 */ assign n138 = n3094;
/* FF 22 10  1 */ always @(posedge n1, posedge n5) if (n5) n1622 <= 1'b0; else if (1'b1) n1622 <= n3095;
/* FF 21 18  1 */ assign n1592 = n3096;
/* FF 12 15  4 */ assign n463 = n3097;
/* FF 18 24  1 */ assign n1270 = n3098;
/* FF 15  7  5 */ assign n738 = n908;
/* FF 20 14  0 */ assign n3099 = n1567;
/* FF 13  8  6 */ assign n545 = n3100;
/* FF 13 19  7 */ assign n395 = n3101;
/* FF 18 23  5 */ always @(posedge n3) if (n881) io_25_33_0 <= 1'b0 ? 1'b0 : n3102;
/* FF 14 18  6 */ always @(posedge n3, posedge n5) if (n5) n185 <= 1'b0; else if (1'b1) n185 <= n3103;
/* FF 11 15  2 */ assign n325 = n3104;
/* FF 14  7  1 */ always @(negedge io_0_6_1, posedge n5) if (n5) n647 <= 1'b0; else if (1'b1) n647 <= n3105;
/* FF 19 12  6 */ assign n1302 = n1435;
/* FF 12 19  3 */ always @(posedge n3, posedge n5) if (n5) n506 <= 1'b0; else if (n620) n506 <= n3106;
/* FF 14 17  0 */ assign n706 = n3107;
/* FF 17 12  4 */ assign n1066 = n3108;
/* FF 17 23  5 */ assign n1142 = n3109;
/* FF 10 15  0 */ assign n219 = n3110;
/* FF 21 19  6 */ always @(posedge n1, posedge n5) if (n5) n1054 <= 1'b0; else if (n8) n1054 <= n3112;
/* FF 13 23  4 */ assign n3113 = n3114;
/* FF 15  9  3 */ always @(posedge n3, posedge n5) if (n5) n552 <= 1'b0; else if (1'b1) n552 <= n3115;
/* FF 12 14  7 */ assign n449 = n3116;
/* FF  6 16  0 */ assign n83 = n3117;
/* FF 20 13  1 */ assign n3118 = n1557;
/* FF 16 23  1 */ always @(posedge n3, posedge n5) if (n5) n1015 <= 1'b0; else if (n1010) n1015 <= n3119;
/* FF 10 17  4 */ always @(posedge n1) if (1'b1) n227 <= n7 ? 1'b0 : n3120;
/* FF 13 20  6 */ assign n627 = n3121;
/* FF 18 13  3 */ assign n3122 = n1314;
/* FF 20 19  0 */ always @(posedge n3, posedge n5) if (n5) n1371 <= 1'b0; else if (n803) n1371 <= n3123;
/* FF 14 13  7 */ always @(posedge n3, posedge n5) if (n5) n450 <= 1'b0; else if (n690) n450 <= n3124;
/* FF 11 12  3 */ always @(posedge n3, posedge n5) if (n5) n42 <= 1'b0; else if (n26) n42 <= n3125;
/* FF 17 19  2 */ assign n3126 = n3127;
/* FF 19 13  1 */ assign n3128 = n1443;
/* FF 22 17  2 */ assign n3129 = n1731;
/* FF 15 24  2 */ always @(posedge n3, posedge n5) if (n5) n884 <= 1'b0; else if (n2) n884 <= n3130;
/* FF 12 18  0 */ always @(posedge n3) if (1'b1) n484 <= n128 ? 1'b0 : n3131;
/* FF 17 13  7 */ assign n1076 = n3132;
/* FF 14 16  3 */ always @(posedge n3, posedge n5) if (n5) n700 <= 1'b0; else if (1'b1) n700 <= n3133;
/* FF 17 16  4 */ assign n3134 = n1213;
/* FF  7  9  6 */ always @(posedge n1, posedge n5) if (n5) n65 <= 1'b1; else if (1'b1) n65 <= n3135;
/* FF 21 20  7 */ always @(posedge n3, posedge n5) if (n5) n1387 <= 1'b0; else if (n270) n1387 <= n3136;
/* FF 13 24  5 */ assign n3137 = n3138;
/* FF 15 14  2 */ assign n359 = n3139;
/* FF 18 17  6 */ assign n1217 = n3140;
/* FF 12 13  6 */ always @(posedge n3, posedge n5) if (n5) n437 <= 1'b0; else if (n573) n437 <= n3141;
/* FF 16 22  2 */ always @(posedge n3) if (n881) io_33_31_0 <= 1'b0 ? 1'b0 : n3142;
/* FF 10 16  7 */ always @(posedge n1) if (1'b1) n237 <= n7 ? 1'b0 : n3143;
/* FF 13 10  4 */ always @(posedge n1, posedge n5) if (n5) n550 <= 1'b0; else if (1'b1) n550 <= n3144;
/* FF 18 12  0 */ always @(posedge n3, posedge n5) if (n5) n1170 <= 1'b0; else if (n1298) n1170 <= n3145;
/* FF 14 12  4 */ assign n3146 = n773;
/* FF 11 13  4 */ always @(posedge n3, posedge n5) if (n5) n301 <= 1'b0; else if (n441) n301 <= n3147;
/* FF 19 10  0 */ always @(posedge n3, posedge n5) if (n5) n1289 <= 1'b0; else if (n580) n1289 <= n3148;
/* FF 22 16  1 */ assign n3149 = n1722;
/* FF 15 25  5 */ always @(posedge n3, posedge n5) if (n5) n885 <= 1'b0; else if (n2) n885 <= n3150;
/* FF 12 17  1 */ always @(posedge n3) if (1'b1) n469 <= n128 ? 1'b0 : n3151;
/* FF 14 19  2 */ always @(posedge n3, posedge n5) if (n5) n516 <= 1'b0; else if (1'b1) n516 <= n3152;
/* FF 17 14  6 */ assign n3153 = n1198;
/* FF 17 17  7 */ assign n1110 = n3154;
/* FF 21 21  4 */ assign n1611 = n3155;
/* FF 15 15  1 */ always @(posedge n3, posedge n5) if (n5) n786 <= 1'b0; else if (n944) n786 <= n3156;
/* FF 11  9  1 */ always @(posedge n1, posedge n5) if (n5) n136 <= 1'b0; else if (1'b1) n136 <= n3157;
/* FF 16 21  3 */ always @(posedge n3, posedge n5) if (n5) n1001 <= 1'b0; else if (n995) n1001 <= n3158;
/* FF 10 19  6 */ always @(posedge n3, posedge n5) if (n5) n253 <= 1'b0; else if (n359) n253 <= n3159;
/* FF 13 11  3 */ always @(posedge io_0_6_1, posedge n5) if (n5) n560 <= 1'b0; else if (1'b1) n560 <= n3160;
/* FF 13 22  4 */ assign n636 = n3161;
/* FF 18 15  1 */ always @(posedge n3, posedge n5) if (n5) n1200 <= 1'b0; else if (n1199) n1200 <= n3162;
/* FF 20 17  2 */ assign n1457 = n3163;
/* FF 14 15  5 */ assign n591 = n798;
/* FF 11 10  5 */ assign io_6_0_1 = n3164;
/* FF 19 11  3 */ always @(posedge n3, posedge n5) if (n5) n1297 <= 1'b0; else if (n1300) n1297 <= n3165;
/* FF 17 15  1 */ assign n1087 = n3166;
/* FF 19 25  0 */ always @(posedge n3, posedge n5) if (n5) n1374 <= 1'b0; else if (n1012) n1374 <= n3167;
/* FF 17 18  6 */ assign n3168 = n3169;
/* FF 22 13  4 */ assign n1640 = n3170;
/* FF 21 22  5 */ assign n1617 = n3171;
/* FF 15 12  0 */ always @(posedge n3, posedge n5) if (n5) n126 <= 1'b0; else if (1'b1) n126 <= n3172;
/* FF 18 19  4 */ assign n1235 = n3173;
/* FF 11 22  0 */ always @(posedge n3, posedge n5) if (n5) n145 <= 1'b0; else if (n273) n145 <= n3174;
/* FF 16 15  5 */ assign n944 = n3175;
/* FF 16 20  4 */ assign n995 = n3176;
/* FF 13 12  2 */ assign n566 = n3177;
/* FF 15 18  3 */ always @(posedge n3, posedge n5) if (n5) n820 <= 1'b0; else if (n826) n820 <= n3178;
/* FF 20 16  5 */ always @(posedge n3, posedge n5) if (n5) n1448 <= 1'b0; else if (n1455) n1448 <= n3179;
/* FF 12 20  3 */ always @(posedge n3, posedge n5) if (n5) n520 <= 1'b1; else if (n538) n520 <= n3180;
/* FF 17 11  6 */ always @(posedge n3, posedge n5) if (n5) n1061 <= 1'b0; else if (n933) n1061 <= n3181;
/* FF 11 11  6 */ always @(posedge n1, posedge n5) if (n5) n295 <= 1'b0; else if (1'b1) n295 <= n3182;
/* FF 23 14  3 */ always @(posedge n3, posedge n5) if (n5) n1716 <= 1'b0; else if (n127) n1716 <= n3183;
/* FF 21 10  0 */ assign n1534 = n1628;
/* FF 12 23  7 */ assign n3184 = n3185;
/* FF 19 22  1 */ always @(posedge n3, posedge n5) if (n5) n1390 <= 1'b0; else if (1'b1) n1390 <= n3186;
/* FF 16 16  1 */ always @(posedge n3, posedge n5) if (n5) n963 <= 1'b0; else if (n799) n963 <= n3187;
/* FF 22 12  7 */ always @(posedge n3, posedge n5) if (n5) n1209 <= 1'b0; else if (n1077) n1209 <= n3188;
/* FF  7 12  5 */ assign n120 = n3189;
/* FF 18 18  3 */ always @(posedge n3, posedge n5) if (n5) n1224 <= 1'b0; else if (n1117) n1224 <= n3190;
/* FF 20 20  2 */ always @(posedge n3, posedge n5) if (n5) n1150 <= 1'b0; else if (n996) n1150 <= n3191;
/* FF 14 10  7 */ always @(posedge n1, posedge n5) if (n5) n664 <= 1'b0; else if (n672) n664 <= n3192;
/* FF 16 14  6 */ assign n127 = n3193;
/* FF  5 17  4 */ always @(posedge n3, posedge n5) if (n5) n48 <= 1'b0; else if (n4) n48 <= n3194;
/* FF 16 19  5 */ always @(posedge n3, posedge n5) if (n5) n990 <= 1'b0; else if (n801) n990 <= n3195;
/* FF 15 19  0 */ always @(posedge n3, posedge n5) if (n5) n836 <= 1'b0; else if (n629) n836 <= n3196;
/* FF 14  9  3 */ assign n3197 = n750;
/* FF 17 20  7 */ assign n1126 = n3198;
/* FF 23 15  0 */ always @(posedge n3, posedge n5) if (n5) n1459 <= 1'b0; else if (n1654) n1459 <= n3199;
/* FF 24 16  0 */ always @(posedge n3, posedge n5) if (n5) n1322 <= 1'b0; else if (n619) n1322 <= n3200;
/* FF 21 16  6 */ assign n3201 = n1666;
/* FF 21 11  7 */ always @(posedge n3, posedge n5) if (n5) n1181 <= 1'b0; else if (n1631) n1181 <= n3202;
/* FF 12 22  4 */ assign n3203 = n3204;
/* FF 19 23  2 */ always @(posedge n3, posedge n5) if (n5) n729 <= 1'b0; else if (1'b1) n729 <= n3205;
/* FF 22 15  6 */ assign n1655 = n3206;
/* FF 18 21  2 */ always @(posedge n3) if (n881) io_33_3_1 <= 1'b0 ? 1'b0 : n3207;
/* FF 20 11  3 */ always @(posedge n3, posedge n5) if (n5) n1426 <= 1'b0; else if (n1199) n1426 <= n3208;
/* FF 11 20  2 */ assign n389 = n3209;
/* FF 16 13  7 */ assign n938 = n3210;
/* FF  5 18  5 */ always @(posedge n3, posedge n5) if (n5) n57 <= 1'b0; else if (n4) n57 <= n3211;
/* FF 16 18  6 */ always @(posedge n3, posedge n5) if (n5) n861 <= 1'b1; else if (n800) n861 <= n3212;
/* FF 10 20  3 */ always @(posedge n3, posedge n5) if (n5) n262 <= 1'b0; else if (n144) n262 <= n3213;
/* FF 15 16  1 */ assign n793 = n3214;
/* FF 21 15  4 */ assign n1573 = n3215;
/* FF 20 25  6 */ always @(posedge n3, posedge n5) if (n5) n1320 <= 1'b0; else if (n1453) n1320 <= n3216;
/* FF 20 22  7 */ assign n272 = n3217;
/* FF 17 24  7 */ assign n3218 = n3219;
/* FF 23 12  1 */ always @(posedge n3) if (n1301) n1565 <= 1'b0 ? 1'b0 : n3220;
/* FF 24 15  1 */ always @(posedge n3, posedge n5) if (n5) n139 <= 1'b0; else if (n958) n139 <= n3221;
/* FF  7 10  6 */ always @(posedge n1, posedge n5) if (n5) n109 <= 1'b0; else if (1'b1) n109 <= n3222;
/* FF 21 17  5 */ always @(posedge n3, posedge n5) if (n5) n1588 <= 1'b0; else if (n1179) n1588 <= n3223;
/* FF 21 12  6 */ always @(posedge n3, posedge n5) if (n5) n1203 <= 1'b0; else if (n1186) n1203 <= n3224;
/* FF 12 21  5 */ assign n535 = n3225;
/* FF 17 10  2 */ always @(posedge n1, posedge n5) if (n5) n414 <= 1'b0; else if (n8) n414 <= n3226;
/* FF 19 20  3 */ always @(posedge n3, posedge n5) if (n5) n1379 <= 1'b0; else if (1'b1) n1379 <= n3227;
/* FF 22 14  1 */ always @(posedge n3, posedge n5) if (n5) n1642 <= 1'b0; else if (n1651) n1642 <= n3228;
/* FF 18 20  1 */ assign n3229 = n1386;
/* FF 20 10  0 */ always @(posedge n1, posedge n5) if (n5) n41 <= 1'b0; else if (1'b1) n41 <= n3230;
/* FF 23 16  7 */ always @(posedge n3, posedge n5) if (n5) n1412 <= 1'b0; else if (n1653) n1412 <= n3231;
/* FF 11 14  4 */ assign n316 = n3232;
/* FF 16 12  0 */ assign n525 = n3233;
/* FF  5 19  2 */ always @(posedge n3, posedge n5) if (n5) n30 <= 1'b0; else if (n4) n30 <= n3234;
/* FF 16 17  7 */ always @(posedge n3, posedge n5) if (n5) n976 <= 1'b0; else if (n702) n976 <= n3235;
/* FF 15 17  6 */ always @(posedge n3, posedge n5) if (n5) n806 <= 1'b0; else if (n609) n806 <= n3236;
/* FF 20 24  1 */ assign n1522 = n3237;
/* FF 12 12  7 */ always @(posedge io_0_6_1, posedge n5) if (n5) n429 <= 1'b0; else if (n563) n429 <= n3238;
/* FF 20 21  6 */ assign n1293 = n3239;
/* FF 17 22  5 */ assign n1134 = n3240;
/* FF 24 14  2 */ always @(posedge n3, posedge n5) if (n5) n1563 <= 1'b0; else if (n467) n1563 <= n3241;
/* FF 22 10  6 */ always @(posedge n1, posedge n5) if (n5) n1626 <= 1'b0; else if (1'b1) n1626 <= n3242;
/* FF 21 18  4 */ assign n1594 = n3243;
/* FF 21 13  5 */ assign n3244 = n1645;
/* FF 12 15  3 */ assign n462 = n3245;
/* FF 19 21  4 */ always @(posedge n3, posedge n5) if (n5) n1287 <= 1'b1; else if (n1145) n1287 <= n3246;
/* FF 10 11  0 */ always @(posedge n1, posedge n5) if (n5) n201 <= 1'b0; else if (n150) n201 <= n3247;
/* FF 15 21  3 */ assign n872 = n3248;
/* FF 18 23  0 */ always @(posedge n3) if (n881) io_19_33_1 <= 1'b0 ? 1'b0 : n3249;
/* FF 23 17  0 */ always @(posedge n3, posedge n5) if (n5) n1726 <= 1'b0; else if (n619) n1726 <= n3250;
/* FF 11 15  7 */ assign n330 = n3251;
/* FF 14  7  4 */ always @(negedge io_0_6_1, posedge n5) if (n5) n650 <= 1'b0; else if (1'b1) n650 <= n3252;
/* FF 11 18  4 */ assign n370 = n3253;
/* FF 16 11  1 */ always @(posedge n3, posedge n5) if (n5) n924 <= 1'b0; else if (n938) n924 <= n3254;
/* FF 15 22  7 */ assign n3255 = n3256;
/* FF 18  9  3 */ always @(posedge n3, posedge n5) if (n5) n1154 <= 1'b0; else if (n215) n1154 <= n3257;
/* FF 12 19  6 */ always @(posedge n3, posedge n5) if (n5) n509 <= 1'b0; else if (n620) n509 <= n3258;
/* FF  6 11  6 */ always @(posedge n1, posedge n5) if (n5) n73 <= 1'b0; else if (1'b1) n73 <= n3259;
/* FF 17 23  2 */ assign n1139 = n3260;
/* FF 19 17  1 */ assign n3261 = n1477;
/* FF 22 21  2 */ always @(posedge n3, posedge n5) if (n5) n1692 <= 1'b0; else if (n1652) n1692 <= n3262;
/* FF 21 19  3 */ assign n3263 = n1682;
/* FF 21 14  4 */ assign n1560 = n3264;
/* FF  9 16  1 */ assign n165 = n3265;
/* FF 12 14  0 */ assign n442 = n3266;
/* FF 14 20  3 */ always @(posedge n3, posedge n5) if (n5) n527 <= 1'b0; else if (1'b1) n527 <= n3268;
/* FF 19 18  5 */ assign n1357 = n3269;
/* FF 10 10  7 */ assign n3270 = n3271;
/* FF 16 23  4 */ always @(posedge n3, posedge n5) if (n5) n1018 <= 1'b0; else if (n1010) n1018 <= n3272;
/* FF 15 10  2 */ always @(posedge n1, posedge n5) if (n5) n554 <= 1'b0; else if (1'b1) n554 <= n3273;
/* FF 20 19  7 */ always @(posedge n3, posedge n5) if (n5) n1115 <= 1'b0; else if (n803) n1115 <= n3274;
/* FF 20  8  6 */ always @(posedge n1, posedge n5) if (n5) n1423 <= 1'b0; else if (n8) n1423 <= n3275;
/* FF 11 12  6 */ always @(posedge n3, posedge n5) if (n5) n140 <= 1'b0; else if (n26) n140 <= n3276;
/* FF 17 19  7 */ assign n3277 = n3278;
/* FF 11 19  7 */ assign n382 = n3279;
/* FF 16 10  2 */ always @(posedge n1, posedge n5) if (n5) n919 <= 1'b0; else if (n672) n919 <= n3280;
/* FF  9 12  3 */ always @(posedge n1, posedge n5) if (n5) n43 <= 1'b0; else if (1'b1) n43 <= n3281;
/* FF 15 24  5 */ always @(posedge n3, posedge n5) if (n5) n889 <= 1'b0; else if (n2) n889 <= n3282;
/* FF 12 18  5 */ always @(posedge n3) if (1'b1) n488 <= n128 ? 1'b0 : n3283;
/* FF 17 16  3 */ assign n1102 = n3284;
/* FF 19 14  0 */ always @(posedge n3, posedge n5) if (n5) n1316 <= 1'b0; else if (n596) n1316 <= n3285;
/* FF 22 20  1 */ assign n1685 = n3286;
/* FF 16 24  2 */ always @(posedge n3, posedge n5) if (n5) n1023 <= 1'b0; else if (n1010) n1023 <= n3287;
/* FF 21 20  2 */ always @(posedge n3, posedge n5) if (n5) n1600 <= 1'b0; else if (n270) n1600 <= n3288;
/* FF 12 13  1 */ always @(posedge n3, posedge n5) if (n5) n432 <= 1'b1; else if (n573) n432 <= n3289;
/* FF 14 23  2 */ always @(posedge n3, posedge n5) if (n5) n31 <= 1'b0; else if (n538) n31 <= n3290;
/* FF 20 12  3 */ always @(posedge n3, posedge n5) if (n5) n1433 <= 1'b0; else if (n1299) n1433 <= n3291;
/* FF 19 19  6 */ always @(posedge n3, posedge n5) if (n5) n1153 <= 1'b0; else if (n985) n1153 <= n3292;
/* FF 10 13  6 */ always @(posedge n1, posedge n5) if (n5) n210 <= 1'b0; else if (n138) n210 <= n3293;
/* FF 15 11  1 */ always @(posedge n1, posedge n5) if (n5) n762 <= 1'b0; else if (1'b1) n762 <= n3294;
/* FF 20 18  4 */ always @(posedge n3, posedge n5) if (n5) n1238 <= 1'b0; else if (n1369) n1238 <= n3295;
/* FF 20 15  7 */ assign n933 = n3296;
/* FF 11 13  1 */ always @(posedge n3, posedge n5) if (n5) n298 <= 1'b0; else if (n441) n298 <= n3297;
/* FF 11 16  6 */ always @(posedge n3, posedge n5) if (n5) n343 <= 1'b0; else if (1'b1) n343 <= n3298;
/* FF 13  7  3 */ assign io_0_6_0 = n3299;
/* FF 15 25  2 */ always @(posedge n3, posedge n5) if (n5) n894 <= 1'b0; else if (n2) n894 <= n3300;
/* FF 18 11  1 */ always @(posedge n3, posedge n5) if (n5) n1160 <= 1'b0; else if (n1179) n1160 <= n3301;
/* FF 15 20  5 */ assign n858 = n3302;
/* FF 12 17  4 */ always @(posedge n3) if (1'b1) n472 <= n128 ? 1'b0 : n3303;
/* FF 17 17  0 */ assign n1105 = n3304;
/* FF 19 15  3 */ assign n3305 = n1464;
/* FF 22 23  0 */ always @(posedge n3, posedge n5) if (n5) n1351 <= 1'b0; else if (n1656) n1351 <= n3306;
/* FF 21 21  1 */ assign n3307 = n1696;
/* FF  9 18  3 */ always @(posedge n3, posedge n5) if (n5) n178 <= 1'b1; else if (n172) n178 <= n3308;
/* FF 14 22  5 */ always @(posedge n3, posedge n5) if (n5) n725 <= 1'b0; else if (n704) n725 <= n3309;
/* FF 11  9  6 */ assign n279 = n408;
/* FF 19 16  7 */ always @(posedge n3, posedge n5) if (n5) n952 <= 1'b0; else if (n949) n952 <= n3310;
/* FF 16 21  6 */ always @(posedge n3, posedge n5) if (n5) n1004 <= 1'b0; else if (n995) n1004 <= n3311;
/* FF 15  8  0 */ assign n3312 = n912;
/* FF 20 17  5 */ always @(posedge n3, posedge n5) if (n5) n1472 <= 1'b0; else if (n793) n1472 <= n3313;
/* FF  6 12  4 */ assign n78 = n123;
/* FF 20 14  4 */ assign n3314 = n1570;
/* FF 23 20  3 */ always @(posedge n3, posedge n5) if (n5) n1506 <= 1'b0; else if (n1655) n1506 <= n3315;
/* FF 11 10  0 */ assign n282 = n412;
/* FF 14 18  2 */ always @(posedge n3, posedge n5) if (n5) n386 <= 1'b0; else if (1'b1) n386 <= n3316;
/* FF 17 18  1 */ assign n3317 = n3318;
/* FF 19 12  2 */ assign n1299 = n3319;
/* FF 21 22  0 */ assign n1616 = n3320;
/* FF 17 12  0 */ always @(posedge n3, posedge n5) if (n5) n1063 <= 1'b0; else if (n619) n1063 <= n3321;
/* FF 14 17  4 */ assign n3322 = n818;
/* FF 11 22  7 */ always @(posedge n3, posedge n5) if (n5) n404 <= 1'b0; else if (n273) n404 <= n3323;
/* FF 10 15  4 */ always @(posedge n1) if (1'b1) n223 <= n7 ? 1'b0 : n3324;
/* FF 16 20  1 */ assign n619 = n3325;
/* FF 15 18  6 */ always @(posedge n3, posedge n5) if (n5) n823 <= 1'b0; else if (n826) n823 <= n3326;
/* FF 13 23  0 */ assign n3327 = n3328;
/* FF 18 14  3 */ assign n1191 = n3329;
/* FF 20 16  2 */ always @(posedge n3, posedge n5) if (n5) n1466 <= 1'b0; else if (n1455) n1466 <= n3330;
/* FF 20 13  5 */ always @(posedge n3, posedge n5) if (n5) n1439 <= 1'b0; else if (n933) n1439 <= n3331;
/* FF 11 11  3 */ always @(posedge n1, posedge n5) if (n5) n286 <= 1'b0; else if (1'b1) n286 <= n3332;
/* FF 22 18  4 */ assign n3333 = n1738;
/* FF 10 17  0 */ always @(posedge n1) if (1'b1) n242 <= n7 ? 1'b0 : n3334;
/* FF  9 15  6 */ assign n163 = n3335;
/* FF 18 13  7 */ assign n1184 = n3336;
/* FF 12 23  2 */ assign n3337 = n3338;
/* FF 14 13  3 */ always @(posedge n3, posedge n5) if (n5) n685 <= 1'b0; else if (n690) n685 <= n3339;
/* FF 19 22  4 */ always @(posedge n3, posedge n5) if (n5) n1393 <= 1'b0; else if (1'b1) n1393 <= n3340;
/* FF 19 13  5 */ assign n3341 = n1445;
/* FF 22 17  6 */ assign n1669 = n3342;
/* FF 16 16  6 */ always @(posedge n3, posedge n5) if (n5) n967 <= 1'b0; else if (n799) n967 <= n3343;
/* FF 15 13  4 */ assign n776 = n947;
/* FF 20 20  7 */ always @(posedge n3, posedge n5) if (n5) n1281 <= 1'b0; else if (n996) n1281 <= n3344;
/* FF 14 16  7 */ always @(posedge n3, posedge n5) if (n5) n701 <= 1'b0; else if (1'b1) n701 <= n3345;
/* FF 17 13  3 */ assign n3346 = n1188;
/* FF 16 19  0 */ always @(posedge n3, posedge n5) if (n5) n878 <= 1'b0; else if (n801) n878 <= n3347;
/* FF  9 11  3 */ assign n153 = n3348;
/* FF 15 19  5 */ always @(posedge n3, posedge n5) if (n5) n840 <= 1'b1; else if (n629) n840 <= n3349;
/* FF 13 24  1 */ assign n3350 = n3351;
/* FF 18 17  2 */ assign n607 = n3352;
/* FF 15 14  6 */ assign n782 = n957;
/* FF 20 23  3 */ always @(posedge n3) if (n688) n1519 <= 1'b0 ? 1'b0 : n3353;
/* FF 10 16  3 */ always @(posedge n1) if (1'b1) n233 <= n7 ? 1'b0 : n3354;
/* FF 13 10  0 */ always @(posedge n1, posedge n5) if (n5) n548 <= 1'b0; else if (1'b1) n548 <= n3355;
/* FF 18 12  4 */ always @(posedge n3, posedge n5) if (n5) n1173 <= 1'b0; else if (n1298) n1173 <= n3356;
/* FF 12 22  1 */ assign n3357 = n3358;
/* FF 14 12  0 */ assign n3359 = n772;
/* FF 19 23  7 */ always @(posedge n3, posedge n5) if (n5) n1148 <= 1'b0; else if (1'b1) n1148 <= n3360;
/* FF 19 10  4 */ always @(posedge n3, posedge n5) if (n5) n1291 <= 1'b0; else if (n580) n1291 <= n3361;
/* FF 22 16  5 */ assign n3362 = n1724;
/* FF 20 11  6 */ always @(posedge n3, posedge n5) if (n5) n1096 <= 1'b0; else if (n1199) n1096 <= n3363;
/* FF 17 14  2 */ always @(posedge n3, posedge n5) if (n5) n1080 <= 1'b0; else if (n958) n1080 <= n3364;
/* FF 14 19  6 */ always @(posedge n3, posedge n5) if (n5) n188 <= 1'b0; else if (1'b1) n188 <= n3365;
/* FF 19 24  3 */ always @(posedge n3, posedge n5) if (n5) n1408 <= 1'b0; else if (n1025) n1408 <= n3366;
/* FF 11 20  5 */ assign n392 = n3367;
/* FF 16 18  3 */ always @(posedge n3, posedge n5) if (n5) n981 <= 1'b1; else if (n800) n981 <= n3368;
/* FF 15 16  4 */ assign n492 = n3369;
/* FF 15 15  5 */ always @(posedge n3, posedge n5) if (n5) n789 <= 1'b0; else if (n944) n789 <= n3370;
/* FF 18 16  1 */ always @(posedge n1, posedge n5) if (n5) n709 <= 1'b0; else if (n8) n709 <= n3371;
/* FF 20 22  0 */ assign n1503 = n3372;
/* FF 17 24  2 */ assign n3373 = n3374;
/* FF 10 19  2 */ always @(posedge n3, posedge n5) if (n5) n249 <= 1'b0; else if (n359) n249 <= n3375;
/* FF 18 15  5 */ assign n3376 = n1335;
/* FF 12 21  0 */ assign n530 = n3377;
/* FF 14 15  1 */ always @(posedge n3) if (n688) n693 <= 1'b0 ? 1'b0 : n3379;
/* FF 19 20  6 */ assign n1012 = n3380;
/* FF 19 11  7 */ always @(posedge n3, posedge n5) if (n5) n940 <= 1'b0; else if (n1300) n940 <= n3381;
/* FF 22 19  4 */ assign n1310 = n3382;
/* FF 24 18  2 */ always @(posedge n1, posedge n5) if (n5) n1219 <= 1'b0; else if (n8) n1219 <= n3383;
/* FF 17 15  5 */ assign n3384 = n1207;
/* FF 16 17  2 */ always @(posedge n3, posedge n5) if (n5) n971 <= 1'b0; else if (n702) n971 <= n3385;
/* FF 22 13  0 */ assign n3386 = n1713;
/* FF 15 17  3 */ always @(posedge n3, posedge n5) if (n5) n811 <= 1'b0; else if (n609) n811 <= n3387;
/* FF 15 12  4 */ assign n768 = n3388;
/* FF 18 19  0 */ assign n1232 = n3389;
/* FF 20 21  1 */ always @(posedge n3, posedge n5) if (n5) n1496 <= 1'b0; else if (n1012) n1496 <= n3390;
/* FF 17 25  1 */ always @(posedge n1, posedge n5) if (n5) n575 <= 1'b0; else if (n8) n575 <= n3391;
/* FF 16 15  1 */ assign n958 = n3392;
/* FF 23 13  3 */ always @(posedge n3, posedge n5) if (n5) n1243 <= 1'b0; else if (n793) n1243 <= n3393;
/* FF 24 14  7 */ always @(posedge n3, posedge n5) if (n5) n695 <= 1'b0; else if (n467) n695 <= n3394;
/* FF 17 11  2 */ assign n1058 = n3395;
/* FF 19 21  1 */ always @(posedge n3, posedge n5) if (n5) n755 <= 1'b1; else if (n1145) n755 <= n3396;
/* FF 11 17  7 */ assign n357 = n3397;
/* FF 23 14  7 */ always @(posedge n3, posedge n5) if (n5) n978 <= 1'b0; else if (n127) n978 <= n3398;
/* FF 24 17  3 */ always @(posedge n3, posedge n5) if (n5) n1226 <= 1'b0; else if (n1454) n1226 <= n3399;
/* FF 17  8  4 */ always @(posedge n3, posedge n5) if (n5) n911 <= 1'b0; else if (1'b1) n911 <= n3400;
/* FF 11 18  3 */ assign n369 = n3401;
/* FF 22 12  3 */ always @(posedge n3, posedge n5) if (n5) n1635 <= 1'b0; else if (n1077) n1635 <= n3402;
/* FF 13 16  5 */ always @(posedge n3, posedge n5) if (n5) n587 <= 1'b0; else if (n492) n587 <= n3403;
/* FF 15 22  2 */ assign n3404 = n3405;
/* FF 18  9  6 */ always @(posedge n3, posedge n5) if (n5) n1158 <= 1'b0; else if (n215) n1158 <= n3406;
/* FF 18 18  7 */ assign n1195 = n3407;
/* FF  6 11  1 */ always @(posedge n1, posedge n5) if (n5) n68 <= 1'b0; else if (1'b1) n68 <= n3408;
/* FF 23 18  1 */ always @(posedge n3, posedge n5) if (n5) n1690 <= 1'b0; else if (n1117) n1690 <= n3409;
/* FF 14 10  3 */ always @(posedge n1, posedge n5) if (n5) n661 <= 1'b0; else if (n672) n661 <= n3410;
/* FF 19 17  6 */ assign n1347 = n3411;
/* FF 16 14  2 */ assign n580 = n3412;
/* FF  5 17  0 */ always @(posedge n3, posedge n5) if (n5) n45 <= 1'b0; else if (n4) n45 <= n3413;
/* FF 14 20  4 */ always @(posedge n3, posedge n5) if (n5) n189 <= 1'b0; else if (1'b1) n189 <= n3414;
/* FF 17 20  3 */ assign n1122 = n3415;
/* FF 19 18  0 */ always @(posedge n3, posedge n5) if (n5) n1355 <= 1'b0; else if (n596) n1355 <= n3416;
/* FF 23 15  4 */ always @(posedge n3, posedge n5) if (n5) n1720 <= 1'b0; else if (n1654) n1720 <= n3417;
/* FF 21 16  2 */ assign n1580 = n3418;
/* FF 18 22  4 */ assign n1145 = n3419;
/* FF 11 19  0 */ assign n375 = n3420;
/* FF 22 15  2 */ assign n1369 = n3421;
/* FF 13 17  6 */ assign n495 = n3422;
/* FF 18 21  6 */ always @(posedge n3) if (n881) io_33_5_0 <= 1'b0 ? 1'b0 : n3423;
/* FF 19 14  7 */ assign n1319 = n3424;
/* FF 16 13  3 */ always @(posedge n3, posedge n5) if (n5) n244 <= 1'b0; else if (n321) n244 <= n3425;
/* FF  5 18  1 */ always @(posedge n3, posedge n5) if (n5) n53 <= 1'b0; else if (n4) n53 <= n3426;
/* FF 10 20  7 */ always @(posedge n3, posedge n5) if (n5) n266 <= 1'b1; else if (n144) n266 <= n3427;
/* FF 13 14  4 */ always @(posedge n3, posedge n5) if (n5) n574 <= 1'b0; else if (n580) n574 <= n3428;
/* FF 21 15  0 */ assign n1571 = n3429;
/* FF 20 25  2 */ always @(posedge n3, posedge n5) if (n5) n1533 <= 1'b0; else if (n1453) n1533 <= n3430;
/* FF 17 21  0 */ assign n1127 = n3431;
/* FF 19 19  3 */ always @(posedge n3, posedge n5) if (n5) n1368 <= 1'b0; else if (n985) n1368 <= n3432;
/* FF 23 12  5 */ always @(posedge n3) if (n1301) n502 <= 1'b0 ? 1'b0 : n3433;
/* FF 21 17  1 */ always @(posedge n3, posedge n5) if (n5) n1585 <= 1'b0; else if (n1179) n1585 <= n3434;
/* FF 18 25  5 */ assign n1278 = n3435;
/* FF 20 15  2 */ assign n1455 = n3436;
/* FF 11 16  1 */ always @(posedge n3, posedge n5) if (n5) n181 <= 1'b0; else if (1'b1) n181 <= n3437;
/* FF 22 14  5 */ always @(posedge n3, posedge n5) if (n5) n1449 <= 1'b0; else if (n1651) n1449 <= n3438;
/* FF 13 18  7 */ assign n384 = n3439;
/* FF 15 20  0 */ assign n853 = n3440;
/* FF 18 20  5 */ assign n1247 = n3442;
/* FF 23 16  3 */ always @(posedge n3, posedge n5) if (n5) n1484 <= 1'b0; else if (n1653) n1484 <= n3443;
/* FF 11 14  0 */ assign n3444 = n3445;
/* FF 16  7  5 */ always @(negedge io_0_6_1, posedge n5) if (n5) n905 <= 1'b0; else if (1'b1) n905 <= n3447;
/* FF 19 15  4 */ assign n1328 = n3448;
/* FF 16 12  4 */ assign n538 = n3449;
/* FF 10 23  6 */ always @(posedge n3, posedge n5) if (n5) n271 <= 1'b0; else if (n273) n271 <= n3450;
/* FF 12 12  3 */ always @(posedge io_0_6_1, posedge n5) if (n5) n426 <= 1'b0; else if (n563) n426 <= n3451;
/* FF 14 22  2 */ always @(posedge n3, posedge n5) if (n5) n723 <= 1'b0; else if (n704) n723 <= n3452;
/* FF 17 22  1 */ assign n1130 = n3453;
/* FF 19 16  2 */ always @(posedge n3, posedge n5) if (n5) n1331 <= 1'b0; else if (n949) n1331 <= n3454;
/* FF 22 10  2 */ always @(posedge n1, posedge n5) if (n5) n1623 <= 1'b0; else if (1'b1) n1623 <= n3455;
/* FF  7 11  1 */ always @(posedge n1, posedge n5) if (n5) n110 <= 1'b0; else if (1'b1) n110 <= n3456;
/* FF 21 18  0 */ assign n3457 = n1673;
/* FF 12 15  7 */ assign n466 = n3458;
/* FF 18 24  6 */ always @(posedge n3, posedge n5) if (n5) n1272 <= 1'b0; else if (n1012) n1272 <= n3459;
/* FF 15  7  2 */ always @(negedge io_0_6_1, posedge n5) if (n5) n735 <= 1'b0; else if (1'b1) n735 <= n3460;
/* FF 20 14  1 */ assign n3461 = n1568;
/* FF 13 19  0 */ assign n267 = n3462;
/* FF 18 23  4 */ always @(posedge n3) if (n881) io_33_28_0 <= 1'b0 ? 1'b0 : n3463;
/* FF 14 18  7 */ always @(posedge n3, posedge n5) if (n5) n184 <= 1'b0; else if (1'b1) n184 <= n3464;
/* FF 23 17  4 */ assign n1728 = n3465;
/* FF 11 15  3 */ assign n326 = n3466;
/* FF 14  7  0 */ always @(negedge io_0_6_1, posedge n5) if (n5) n646 <= 1'b0; else if (1'b1) n646 <= n3467;
/* FF 19 12  5 */ assign n1077 = n3469;
/* FF 16 11  5 */ always @(posedge n3, posedge n5) if (n5) n926 <= 1'b0; else if (n938) n926 <= n3470;
/* FF 12 19  2 */ always @(posedge n3, posedge n5) if (n5) n505 <= 1'b0; else if (n620) n505 <= n3471;
/* FF 17 12  7 */ assign n1069 = n3472;
/* FF 14 17  3 */ assign n3473 = n817;
/* FF 17 23  6 */ assign n1143 = n3474;
/* FF 13 23  5 */ assign n3475 = n3476;
/* FF 12 14  4 */ assign n446 = n3477;
/* FF 20 13  0 */ assign n1436 = n3478;
/* FF 16 23  0 */ always @(posedge n3, posedge n5) if (n5) n1014 <= 1'b0; else if (n1010) n1014 <= n3479;
/* FF 10 17  7 */ assign n3480 = n3481;
/* FF 13 20  1 */ assign n622 = n3482;
/* FF 18 13  2 */ assign n3483 = n1313;
/* FF 20 19  3 */ always @(posedge n3, posedge n5) if (n5) n1249 <= 1'b0; else if (n803) n1249 <= n3484;
/* FF 14 13  6 */ always @(posedge n3, posedge n5) if (n5) n677 <= 1'b0; else if (n690) n677 <= n3485;
/* FF 23 22  5 */ always @(posedge n3, posedge n5) if (n5) n1035 <= 1'b0; else if (n793) n1035 <= n3486;
/* FF 17 19  3 */ assign n3487 = n3488;
/* FF 19 13  2 */ assign n3489 = n1444;
/* FF 16 10  6 */ always @(posedge n1, posedge n5) if (n5) n922 <= 1'b0; else if (n672) n922 <= n3490;
/* FF 15 24  1 */ always @(posedge n3, posedge n5) if (n5) n883 <= 1'b0; else if (n2) n883 <= n3491;
/* FF 12 18  1 */ always @(posedge n3) if (1'b1) n485 <= n128 ? 1'b0 : n3492;
/* FF 14 16  0 */ assign n697 = n3493;
/* FF 17 13  4 */ assign n794 = n3494;
/* FF 21 20  6 */ always @(posedge n3, posedge n5) if (n5) n1607 <= 1'b0; else if (n270) n1607 <= n3495;
/* FF 13 24  4 */ assign n3496 = n3497;
/* FF  9 17  6 */ always @(posedge n3, posedge n5) if (n5) n129 <= 1'b0; else if (n172) n129 <= n3498;
/* FF 12 13  5 */ always @(posedge n3, posedge n5) if (n5) n436 <= 1'b0; else if (n573) n436 <= n3499;
/* FF 18 26  0 */ assign n2 = n3500;
/* FF 16 22  3 */ assign n4 = n3501;
/* FF 10 16  4 */ always @(posedge n1) if (1'b1) n234 <= n7 ? 1'b0 : n3502;
/* FF 18 12  1 */ always @(posedge n3, posedge n5) if (n5) n1171 <= 1'b0; else if (n1298) n1171 <= n3503;
/* FF  6 13  3 */ assign n81 = n3504;
/* FF 20 18  0 */ assign n1093 = n3505;
/* FF 14 12  5 */ assign n3506 = n774;
/* FF 11 13  5 */ always @(posedge n3, posedge n5) if (n5) n302 <= 1'b0; else if (n441) n302 <= n3507;
/* FF 15 25  6 */ always @(posedge n3, posedge n5) if (n5) n896 <= 1'b0; else if (n2) n896 <= n3508;
/* FF 12 17  0 */ always @(posedge n3) if (1'b1) n468 <= n128 ? 1'b0 : n3509;
/* FF 17 14  5 */ always @(posedge n3, posedge n5) if (n5) n1082 <= 1'b0; else if (n958) n1082 <= n3511;
/* FF 14 19  1 */ always @(posedge n3, posedge n5) if (n5) n268 <= 1'b0; else if (1'b1) n268 <= n3512;
/* FF 17 17  4 */ always @(posedge n3, posedge n5) if (n5) n1108 <= 1'b0; else if (n985) n1108 <= n3513;
/* FF 21 21  5 */ assign n1612 = n3514;
/* FF 16 21  2 */ always @(posedge n3, posedge n5) if (n5) n1000 <= 1'b0; else if (n995) n1000 <= n3515;
/* FF 10 19  5 */ always @(posedge n3, posedge n5) if (n5) n252 <= 1'b0; else if (n359) n252 <= n3516;
/* FF 13 22  3 */ assign n635 = n3517;
/* FF 18 15  0 */ assign n1199 = n3518;
/* FF  6 12  0 */ assign n66 = n3519;
/* FF 20 17  1 */ always @(posedge n3, posedge n5) if (n5) n1469 <= 1'b0; else if (n793) n1469 <= n3520;
/* FF 14 15  4 */ always @(posedge n3) if (n688) n694 <= 1'b0 ? 1'b0 : n3521;
/* FF 23 20  7 */ always @(posedge n3, posedge n5) if (n5) n1262 <= 1'b0; else if (n1655) n1262 <= n3522;
/* FF 19 11  0 */ always @(posedge n3, posedge n5) if (n5) n986 <= 1'b0; else if (n1300) n986 <= n3523;
/* FF 17 15  2 */ always @(posedge n3, posedge n5) if (n5) n1088 <= 1'b0; else if (n805) n1088 <= n3524;
/* FF 19 25  1 */ always @(posedge n3, posedge n5) if (n5) n1375 <= 1'b0; else if (n1012) n1375 <= n3525;
/* FF 17 18  5 */ assign n3526 = n3527;
/* FF 22 13  7 */ assign n1456 = n3528;
/* FF 11 22  3 */ always @(posedge n3, posedge n5) if (n5) n401 <= 1'b0; else if (n273) n401 <= n3529;
/* FF 16 15  4 */ assign n803 = n3530;
/* FF 16 20  5 */ assign n629 = n3531;
/* FF 15 18  2 */ always @(posedge n3, posedge n5) if (n5) n819 <= 1'b0; else if (n826) n819 <= n3532;
/* FF 20 16  6 */ always @(posedge n3, posedge n5) if (n5) n1085 <= 1'b0; else if (n1455) n1085 <= n3533;
/* FF 17 11  7 */ always @(posedge n3, posedge n5) if (n5) n1062 <= 1'b0; else if (n933) n1062 <= n3534;
/* FF 11 11  7 */ always @(posedge n1, posedge n5) if (n5) n296 <= 1'b0; else if (1'b1) n296 <= n3535;
/* FF 23 14  2 */ always @(posedge n3, posedge n5) if (n5) n1460 <= 1'b0; else if (n127) n1460 <= n3536;
/* FF 22 18  0 */ assign n3537 = n1736;
/* FF 21 10  7 */ assign n1539 = n3538;
/* FF 12 23  6 */ assign n3539 = n3540;
/* FF 19 22  0 */ always @(posedge n3, posedge n5) if (n5) n1389 <= 1'b0; else if (1'b1) n1389 <= n3541;

endmodule

